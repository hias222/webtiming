<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SG Fürth" version="11.61084">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Nürnberg" name="Bayerische Kurzbahnmeisterschaften 2016" course="SCM" deadline="2016-10-26" hostclub="SG Mittelfranken" organizer="Bayerischer Schwimmverband e.V." organizer.url="http://www.bayerischer-schwimmverband.de/schwimmen" reservecount="4" startmethod="1" timing="AUTOMATIC" nation="GER">
      <AGEDATE value="2016-11-06" type="YEAR" />
      <POOL name="90471 Nürnberg, Hallenbad Langwasser, Breslauer Str. 251, Eingang Gleiwitzer Straße" lanemin="1" lanemax="6" />
      <FACILITY city="Nürnberg" name="90471 Nürnberg, Hallenbad Langwasser, Breslauer Str. 251, Eingang Gleiwitzer Straße" nation="GER" />
      <POINTTABLE pointtableid="3009" name="FINA Point Scoring" version="2016" />
      <CONTACT city="Fürth" email="meldungen@sgfuerth.de" name="Matthias Fuchs" phone="09118101172" street="Lavendelweg 47" zip="90768" />
      <QUALIFY from="2016-01-01" until="2016-10-28" />
      <SESSIONS>
        <SESSION date="2016-11-05" daytime="10:00" number="1" officialmeeting="09:30" teamleadermeeting="09:30" warmupfrom="08:30" warmupuntil="09:50">
          <EVENTS>
            <EVENT eventid="1841" daytime="14:05" gender="F" number="15" order="26" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1842" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3504" />
                    <RANKING order="2" place="2" resultid="3023" />
                    <RANKING order="3" place="3" resultid="3834" />
                    <RANKING order="4" place="4" resultid="3061" />
                    <RANKING order="5" place="5" resultid="2925" />
                    <RANKING order="6" place="6" resultid="2948" />
                    <RANKING order="7" place="7" resultid="3301" />
                    <RANKING order="8" place="8" resultid="3978" />
                    <RANKING order="9" place="9" resultid="3605" />
                    <RANKING order="10" place="10" resultid="3295" />
                    <RANKING order="11" place="11" resultid="3965" />
                    <RANKING order="12" place="12" resultid="2479" />
                    <RANKING order="13" place="13" resultid="3960" />
                    <RANKING order="14" place="14" resultid="3043" />
                    <RANKING order="15" place="15" resultid="3861" />
                    <RANKING order="16" place="16" resultid="4145" />
                    <RANKING order="17" place="17" resultid="2601" />
                    <RANKING order="18" place="18" resultid="4606" />
                    <RANKING order="19" place="19" resultid="3953" />
                    <RANKING order="20" place="20" resultid="2564" />
                    <RANKING order="21" place="21" resultid="3006" />
                    <RANKING order="22" place="22" resultid="2614" />
                    <RANKING order="23" place="23" resultid="2792" />
                    <RANKING order="24" place="24" resultid="4045" />
                    <RANKING order="25" place="25" resultid="3923" />
                    <RANKING order="26" place="26" resultid="3617" />
                    <RANKING order="27" place="27" resultid="3415" />
                    <RANKING order="28" place="28" resultid="4598" />
                    <RANKING order="29" place="29" resultid="3388" />
                    <RANKING order="30" place="30" resultid="3769" />
                    <RANKING order="31" place="31" resultid="4073" />
                    <RANKING order="32" place="32" resultid="4006" />
                    <RANKING order="33" place="33" resultid="2988" />
                    <RANKING order="34" place="34" resultid="3844" />
                    <RANKING order="35" place="-1" resultid="2816" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4779" daytime="14:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4780" daytime="14:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4781" daytime="14:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4782" daytime="14:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4783" daytime="14:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4784" daytime="14:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1763" daytime="10:50" gender="M" number="4" order="7" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1764" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3597" />
                    <RANKING order="2" place="2" resultid="4115" />
                    <RANKING order="3" place="3" resultid="3128" />
                    <RANKING order="4" place="4" resultid="3525" />
                    <RANKING order="5" place="5" resultid="2810" />
                    <RANKING order="6" place="6" resultid="3508" />
                    <RANKING order="7" place="7" resultid="3010" />
                    <RANKING order="8" place="8" resultid="3319" />
                    <RANKING order="9" place="9" resultid="2431" />
                    <RANKING order="10" place="10" resultid="2631" />
                    <RANKING order="11" place="11" resultid="3940" />
                    <RANKING order="12" place="12" resultid="3028" />
                    <RANKING order="13" place="13" resultid="3760" />
                    <RANKING order="14" place="14" resultid="2462" />
                    <RANKING order="15" place="15" resultid="3675" />
                    <RANKING order="16" place="16" resultid="3932" />
                    <RANKING order="17" place="17" resultid="3826" />
                    <RANKING order="18" place="18" resultid="4610" />
                    <RANKING order="19" place="19" resultid="2757" />
                    <RANKING order="20" place="20" resultid="4131" />
                    <RANKING order="21" place="21" resultid="3558" />
                    <RANKING order="22" place="22" resultid="2547" />
                    <RANKING order="23" place="23" resultid="3671" />
                    <RANKING order="24" place="24" resultid="4020" />
                    <RANKING order="25" place="25" resultid="2413" />
                    <RANKING order="26" place="26" resultid="4125" />
                    <RANKING order="27" place="27" resultid="2897" />
                    <RANKING order="28" place="28" resultid="2821" />
                    <RANKING order="29" place="29" resultid="3449" />
                    <RANKING order="30" place="30" resultid="3288" />
                    <RANKING order="31" place="31" resultid="3850" />
                    <RANKING order="32" place="32" resultid="2400" />
                    <RANKING order="33" place="33" resultid="3471" />
                    <RANKING order="34" place="34" resultid="3657" />
                    <RANKING order="35" place="35" resultid="2408" />
                    <RANKING order="36" place="36" resultid="3403" />
                    <RANKING order="37" place="37" resultid="2779" />
                    <RANKING order="38" place="38" resultid="4575" />
                    <RANKING order="39" place="39" resultid="2439" />
                    <RANKING order="40" place="40" resultid="3970" />
                    <RANKING order="41" place="41" resultid="3485" />
                    <RANKING order="42" place="42" resultid="3742" />
                    <RANKING order="43" place="43" resultid="2738" />
                    <RANKING order="44" place="44" resultid="2514" />
                    <RANKING order="45" place="45" resultid="3747" />
                    <RANKING order="46" place="46" resultid="3898" />
                    <RANKING order="47" place="-1" resultid="2639" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4696" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4697" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4698" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4699" daytime="10:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4700" daytime="10:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4701" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4702" daytime="11:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4703" daytime="11:00" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1813" daytime="12:45" gender="F" number="11" order="19" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1814" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3532" />
                    <RANKING order="2" place="2" resultid="3927" />
                    <RANKING order="3" place="3" resultid="4080" />
                    <RANKING order="4" place="4" resultid="4075" />
                    <RANKING order="5" place="5" resultid="2941" />
                    <RANKING order="6" place="6" resultid="2498" />
                    <RANKING order="7" place="7" resultid="4167" />
                    <RANKING order="8" place="8" resultid="2456" />
                    <RANKING order="9" place="9" resultid="2962" />
                    <RANKING order="10" place="10" resultid="4621" />
                    <RANKING order="11" place="11" resultid="3015" />
                    <RANKING order="12" place="12" resultid="2701" />
                    <RANKING order="13" place="13" resultid="4955" />
                    <RANKING order="14" place="-1" resultid="3576" />
                    <RANKING order="15" place="-1" resultid="3877" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4745" daytime="12:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4746" daytime="12:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4747" daytime="12:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1792" daytime="11:50" gender="M" number="8" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1793" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3628" />
                    <RANKING order="2" place="2" resultid="2979" />
                    <RANKING order="3" place="3" resultid="3166" />
                    <RANKING order="4" place="4" resultid="2569" />
                    <RANKING order="5" place="5" resultid="2929" />
                    <RANKING order="6" place="6" resultid="3520" />
                    <RANKING order="7" place="7" resultid="3053" />
                    <RANKING order="8" place="8" resultid="2731" />
                    <RANKING order="9" place="9" resultid="3818" />
                    <RANKING order="10" place="10" resultid="3775" />
                    <RANKING order="11" place="11" resultid="4637" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4726" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4727" daytime="12:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1827" daytime="13:15" gender="F" number="13" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1828" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3587" />
                    <RANKING order="2" place="2" resultid="3109" />
                    <RANKING order="3" place="3" resultid="2942" />
                    <RANKING order="4" place="4" resultid="2499" />
                    <RANKING order="5" place="5" resultid="3581" />
                    <RANKING order="6" place="6" resultid="3610" />
                    <RANKING order="7" place="7" resultid="4195" />
                    <RANKING order="8" place="8" resultid="3548" />
                    <RANKING order="9" place="9" resultid="3538" />
                    <RANKING order="10" place="10" resultid="3754" />
                    <RANKING order="11" place="11" resultid="4067" />
                    <RANKING order="12" place="12" resultid="3204" />
                    <RANKING order="13" place="13" resultid="2885" />
                    <RANKING order="14" place="14" resultid="3837" />
                    <RANKING order="15" place="15" resultid="4201" />
                    <RANKING order="16" place="16" resultid="4229" />
                    <RANKING order="17" place="17" resultid="3334" />
                    <RANKING order="18" place="18" resultid="3177" />
                    <RANKING order="19" place="19" resultid="3048" />
                    <RANKING order="20" place="20" resultid="3736" />
                    <RANKING order="21" place="21" resultid="2563" />
                    <RANKING order="22" place="22" resultid="3922" />
                    <RANKING order="23" place="23" resultid="2691" />
                    <RANKING order="24" place="24" resultid="3720" />
                    <RANKING order="25" place="25" resultid="2934" />
                    <RANKING order="26" place="26" resultid="4136" />
                    <RANKING order="27" place="27" resultid="3383" />
                    <RANKING order="28" place="28" resultid="2866" />
                    <RANKING order="29" place="29" resultid="3811" />
                    <RANKING order="30" place="30" resultid="3257" />
                    <RANKING order="31" place="31" resultid="2509" />
                    <RANKING order="32" place="32" resultid="4622" />
                    <RANKING order="33" place="33" resultid="3396" />
                    <RANKING order="34" place="34" resultid="3069" />
                    <RANKING order="35" place="35" resultid="2724" />
                    <RANKING order="36" place="36" resultid="4262" />
                    <RANKING order="37" place="37" resultid="3242" />
                    <RANKING order="38" place="-1" resultid="2577" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4758" daytime="13:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4759" daytime="13:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4760" daytime="13:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4761" daytime="13:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4762" daytime="13:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4763" daytime="13:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4764" daytime="13:50" number="7" order="7" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1820" daytime="12:55" gender="M" number="12" order="20" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1821" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3074" />
                    <RANKING order="2" place="2" resultid="3509" />
                    <RANKING order="3" place="3" resultid="3129" />
                    <RANKING order="4" place="4" resultid="3515" />
                    <RANKING order="5" place="5" resultid="3570" />
                    <RANKING order="6" place="6" resultid="2464" />
                    <RANKING order="7" place="7" resultid="3761" />
                    <RANKING order="8" place="8" resultid="3665" />
                    <RANKING order="9" place="9" resultid="4593" />
                    <RANKING order="10" place="10" resultid="3998" />
                    <RANKING order="11" place="11" resultid="3088" />
                    <RANKING order="12" place="12" resultid="2853" />
                    <RANKING order="13" place="13" resultid="3189" />
                    <RANKING order="14" place="14" resultid="2415" />
                    <RANKING order="15" place="15" resultid="2606" />
                    <RANKING order="16" place="16" resultid="3934" />
                    <RANKING order="17" place="17" resultid="3554" />
                    <RANKING order="18" place="18" resultid="4612" />
                    <RANKING order="19" place="19" resultid="2967" />
                    <RANKING order="20" place="20" resultid="3559" />
                    <RANKING order="21" place="21" resultid="2570" />
                    <RANKING order="22" place="22" resultid="3377" />
                    <RANKING order="23" place="23" resultid="3941" />
                    <RANKING order="24" place="24" resultid="3095" />
                    <RANKING order="25" place="25" resultid="3167" />
                    <RANKING order="26" place="26" resultid="2774" />
                    <RANKING order="27" place="27" resultid="2780" />
                    <RANKING order="28" place="28" resultid="2830" />
                    <RANKING order="29" place="29" resultid="2549" />
                    <RANKING order="30" place="30" resultid="3409" />
                    <RANKING order="31" place="31" resultid="3971" />
                    <RANKING order="32" place="32" resultid="3889" />
                    <RANKING order="33" place="33" resultid="2653" />
                    <RANKING order="34" place="34" resultid="3489" />
                    <RANKING order="35" place="35" resultid="4029" />
                    <RANKING order="36" place="36" resultid="3827" />
                    <RANKING order="37" place="37" resultid="3852" />
                    <RANKING order="38" place="38" resultid="4126" />
                    <RANKING order="39" place="39" resultid="3404" />
                    <RANKING order="40" place="40" resultid="2930" />
                    <RANKING order="41" place="41" resultid="2646" />
                    <RANKING order="42" place="42" resultid="4190" />
                    <RANKING order="43" place="43" resultid="3819" />
                    <RANKING order="44" place="44" resultid="2515" />
                    <RANKING order="45" place="-1" resultid="2640" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4749" daytime="12:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4750" daytime="13:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4751" daytime="13:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4752" daytime="13:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4753" daytime="13:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4754" daytime="13:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4755" daytime="13:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4756" daytime="13:15" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1756" daytime="10:40" gender="F" number="3" order="5" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1757" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3141" />
                    <RANKING order="2" place="2" resultid="3022" />
                    <RANKING order="3" place="3" resultid="2947" />
                    <RANKING order="4" place="4" resultid="4166" />
                    <RANKING order="5" place="5" resultid="4025" />
                    <RANKING order="6" place="6" resultid="3294" />
                    <RANKING order="7" place="7" resultid="2924" />
                    <RANKING order="8" place="8" resultid="3832" />
                    <RANKING order="9" place="9" resultid="2477" />
                    <RANKING order="10" place="10" resultid="3299" />
                    <RANKING order="11" place="11" resultid="4256" />
                    <RANKING order="12" place="12" resultid="3436" />
                    <RANKING order="13" place="13" resultid="2814" />
                    <RANKING order="14" place="14" resultid="4150" />
                    <RANKING order="15" place="15" resultid="3951" />
                    <RANKING order="16" place="16" resultid="4042" />
                    <RANKING order="17" place="17" resultid="3413" />
                    <RANKING order="18" place="18" resultid="2561" />
                    <RANKING order="19" place="19" resultid="3429" />
                    <RANKING order="20" place="20" resultid="3859" />
                    <RANKING order="21" place="21" resultid="3040" />
                    <RANKING order="22" place="22" resultid="2600" />
                    <RANKING order="23" place="23" resultid="2613" />
                    <RANKING order="24" place="24" resultid="3425" />
                    <RANKING order="25" place="25" resultid="3959" />
                    <RANKING order="26" place="26" resultid="2472" />
                    <RANKING order="27" place="27" resultid="2762" />
                    <RANKING order="28" place="28" resultid="3767" />
                    <RANKING order="29" place="29" resultid="2485" />
                    <RANKING order="30" place="30" resultid="4144" />
                    <RANKING order="31" place="31" resultid="4605" />
                    <RANKING order="32" place="32" resultid="3616" />
                    <RANKING order="33" place="33" resultid="2589" />
                    <RANKING order="34" place="34" resultid="3695" />
                    <RANKING order="35" place="35" resultid="2791" />
                    <RANKING order="36" place="36" resultid="2803" />
                    <RANKING order="37" place="37" resultid="4072" />
                    <RANKING order="38" place="38" resultid="4596" />
                    <RANKING order="39" place="39" resultid="2987" />
                    <RANKING order="40" place="40" resultid="2592" />
                    <RANKING order="41" place="41" resultid="3921" />
                    <RANKING order="42" place="42" resultid="3004" />
                    <RANKING order="43" place="43" resultid="2767" />
                    <RANKING order="44" place="44" resultid="3843" />
                    <RANKING order="45" place="45" resultid="2506" />
                    <RANKING order="46" place="46" resultid="2714" />
                    <RANKING order="47" place="47" resultid="2520" />
                    <RANKING order="48" place="-1" resultid="3875" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4687" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4688" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4689" daytime="10:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4690" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4691" daytime="10:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4692" daytime="10:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4693" daytime="10:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4694" daytime="10:45" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1785" daytime="11:40" gender="F" number="7" order="13" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1786" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3108" />
                    <RANKING order="2" place="2" resultid="4066" />
                    <RANKING order="3" place="3" resultid="3946" />
                    <RANKING order="4" place="4" resultid="2992" />
                    <RANKING order="5" place="5" resultid="4058" />
                    <RANKING order="6" place="6" resultid="3060" />
                    <RANKING order="7" place="7" resultid="3802" />
                    <RANKING order="8" place="8" resultid="3014" />
                    <RANKING order="9" place="9" resultid="3203" />
                    <RANKING order="10" place="10" resultid="2497" />
                    <RANKING order="11" place="11" resultid="4650" />
                    <RANKING order="12" place="12" resultid="3266" />
                    <RANKING order="13" place="13" resultid="3480" />
                    <RANKING order="14" place="14" resultid="3354" />
                    <RANKING order="15" place="15" resultid="3150" />
                    <RANKING order="16" place="16" resultid="3142" />
                    <RANKING order="17" place="17" resultid="4012" />
                    <RANKING order="18" place="18" resultid="3753" />
                    <RANKING order="19" place="19" resultid="2541" />
                    <RANKING order="20" place="20" resultid="4151" />
                    <RANKING order="21" place="21" resultid="2787" />
                    <RANKING order="22" place="22" resultid="2884" />
                    <RANKING order="23" place="23" resultid="4617" />
                    <RANKING order="24" place="24" resultid="3913" />
                    <RANKING order="25" place="25" resultid="2690" />
                    <RANKING order="26" place="26" resultid="2745" />
                    <RANKING order="27" place="27" resultid="4052" />
                    <RANKING order="28" place="28" resultid="3768" />
                    <RANKING order="29" place="29" resultid="3219" />
                    <RANKING order="30" place="30" resultid="4043" />
                    <RANKING order="31" place="31" resultid="3810" />
                    <RANKING order="32" place="32" resultid="2447" />
                    <RANKING order="33" place="33" resultid="3183" />
                    <RANKING order="34" place="34" resultid="2715" />
                    <RANKING order="35" place="35" resultid="3116" />
                    <RANKING order="36" place="36" resultid="4579" />
                    <RANKING order="37" place="37" resultid="2507" />
                    <RANKING order="38" place="38" resultid="2528" />
                    <RANKING order="39" place="39" resultid="3226" />
                    <RANKING order="40" place="-1" resultid="3032" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4718" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4719" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4720" daytime="11:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4721" daytime="11:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4722" daytime="11:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4723" daytime="11:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4724" daytime="11:45" number="7" order="7" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1749" daytime="10:20" gender="M" number="2" order="3" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1750" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3073" />
                    <RANKING order="2" place="2" resultid="3997" />
                    <RANKING order="3" place="3" resultid="3622" />
                    <RANKING order="4" place="4" resultid="3087" />
                    <RANKING order="5" place="5" resultid="3569" />
                    <RANKING order="6" place="6" resultid="2859" />
                    <RANKING order="7" place="7" resultid="3553" />
                    <RANKING order="8" place="8" resultid="3514" />
                    <RANKING order="9" place="9" resultid="3194" />
                    <RANKING order="10" place="10" resultid="3465" />
                    <RANKING order="11" place="11" resultid="3080" />
                    <RANKING order="12" place="12" resultid="2623" />
                    <RANKING order="13" place="13" resultid="4213" />
                    <RANKING order="14" place="14" resultid="2852" />
                    <RANKING order="15" place="15" resultid="2978" />
                    <RANKING order="16" place="16" resultid="2568" />
                    <RANKING order="17" place="17" resultid="3164" />
                    <RANKING order="18" place="18" resultid="3691" />
                    <RANKING order="19" place="19" resultid="3982" />
                    <RANKING order="20" place="20" resultid="3661" />
                    <RANKING order="21" place="21" resultid="2604" />
                    <RANKING order="22" place="22" resultid="3408" />
                    <RANKING order="23" place="23" resultid="2730" />
                    <RANKING order="24" place="24" resultid="2438" />
                    <RANKING order="25" place="25" resultid="3093" />
                    <RANKING order="26" place="26" resultid="2891" />
                    <RANKING order="27" place="27" resultid="3866" />
                    <RANKING order="28" place="28" resultid="3155" />
                    <RANKING order="29" place="29" resultid="2828" />
                    <RANKING order="30" place="30" resultid="3323" />
                    <RANKING order="31" place="31" resultid="2773" />
                    <RANKING order="32" place="32" resultid="3135" />
                    <RANKING order="33" place="33" resultid="4118" />
                    <RANKING order="34" place="34" resultid="3100" />
                    <RANKING order="35" place="35" resultid="2996" />
                    <RANKING order="36" place="36" resultid="2652" />
                    <RANKING order="37" place="37" resultid="3774" />
                    <RANKING order="38" place="38" resultid="3882" />
                    <RANKING order="39" place="39" resultid="4027" />
                    <RANKING order="40" place="40" resultid="3460" />
                    <RANKING order="41" place="41" resultid="4174" />
                    <RANKING order="42" place="42" resultid="4586" />
                    <RANKING order="43" place="43" resultid="3817" />
                    <RANKING order="44" place="44" resultid="2423" />
                    <RANKING order="45" place="45" resultid="2952" />
                    <RANKING order="46" place="46" resultid="4574" />
                    <RANKING order="47" place="47" resultid="2645" />
                    <RANKING order="48" place="48" resultid="2660" />
                    <RANKING order="49" place="49" resultid="3713" />
                    <RANKING order="50" place="50" resultid="3360" />
                    <RANKING order="51" place="51" resultid="4950" />
                    <RANKING order="52" place="52" resultid="3687" />
                    <RANKING order="53" place="53" resultid="4189" />
                    <RANKING order="54" place="54" resultid="2683" />
                    <RANKING order="55" place="55" resultid="4646" />
                    <RANKING order="56" place="-1" resultid="2638" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4676" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4677" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4678" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4679" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4680" daytime="10:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4681" daytime="10:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4682" daytime="10:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4683" daytime="10:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4684" daytime="10:35" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4685" daytime="10:40" number="10" order="10" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1806" daytime="12:40" gender="M" number="10" order="18" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1807" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3037" />
                    <RANKING order="2" place="2" resultid="3442" />
                    <RANKING order="3" place="3" resultid="2450" />
                    <RANKING order="4" place="4" resultid="4182" />
                    <RANKING order="5" place="5" resultid="3347" />
                    <RANKING order="6" place="6" resultid="2625" />
                    <RANKING order="7" place="7" resultid="4235" />
                    <RANKING order="8" place="8" resultid="3475" />
                    <RANKING order="9" place="9" resultid="3498" />
                    <RANKING order="10" place="10" resultid="3136" />
                    <RANKING order="11" place="11" resultid="2605" />
                    <RANKING order="12" place="12" resultid="3933" />
                    <RANKING order="13" place="13" resultid="3697" />
                    <RANKING order="14" place="14" resultid="2432" />
                    <RANKING order="15" place="15" resultid="3902" />
                    <RANKING order="16" place="16" resultid="2555" />
                    <RANKING order="17" place="17" resultid="2632" />
                    <RANKING order="18" place="18" resultid="2822" />
                    <RANKING order="19" place="19" resultid="2841" />
                    <RANKING order="20" place="20" resultid="3364" />
                    <RANKING order="21" place="21" resultid="3157" />
                    <RANKING order="22" place="22" resultid="3851" />
                    <RANKING order="23" place="23" resultid="2536" />
                    <RANKING order="24" place="24" resultid="4175" />
                    <RANKING order="25" place="25" resultid="2705" />
                    <RANKING order="26" place="26" resultid="2837" />
                    <RANKING order="27" place="27" resultid="2806" />
                    <RANKING order="28" place="28" resultid="3731" />
                    <RANKING order="29" place="29" resultid="3776" />
                    <RANKING order="30" place="30" resultid="2425" />
                    <RANKING order="31" place="31" resultid="2483" />
                    <RANKING order="32" place="32" resultid="2492" />
                    <RANKING order="33" place="33" resultid="2583" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4738" daytime="12:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4739" daytime="12:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4740" daytime="12:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4741" daytime="12:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4742" daytime="12:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4743" daytime="12:45" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1778" daytime="11:25" gender="M" number="6" order="11" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1779" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3563" />
                    <RANKING order="2" place="2" resultid="3466" />
                    <RANKING order="3" place="3" resultid="2624" />
                    <RANKING order="4" place="4" resultid="2860" />
                    <RANKING order="5" place="5" resultid="2463" />
                    <RANKING order="6" place="6" resultid="3664" />
                    <RANKING order="7" place="7" resultid="3094" />
                    <RANKING order="8" place="8" resultid="3441" />
                    <RANKING order="9" place="9" resultid="2997" />
                    <RANKING order="10" place="10" resultid="4234" />
                    <RANKING order="11" place="11" resultid="3313" />
                    <RANKING order="12" place="12" resultid="4214" />
                    <RANKING order="13" place="12" resultid="4592" />
                    <RANKING order="14" place="14" resultid="3276" />
                    <RANKING order="15" place="15" resultid="3993" />
                    <RANKING order="16" place="16" resultid="2414" />
                    <RANKING order="17" place="17" resultid="3165" />
                    <RANKING order="18" place="18" resultid="3081" />
                    <RANKING order="19" place="19" resultid="2847" />
                    <RANKING order="20" place="20" resultid="4138" />
                    <RANKING order="21" place="21" resultid="3346" />
                    <RANKING order="22" place="22" resultid="3461" />
                    <RANKING order="23" place="23" resultid="2440" />
                    <RANKING order="24" place="23" resultid="3376" />
                    <RANKING order="25" place="25" resultid="3730" />
                    <RANKING order="26" place="26" resultid="2548" />
                    <RANKING order="27" place="27" resultid="3901" />
                    <RANKING order="28" place="28" resultid="2953" />
                    <RANKING order="29" place="29" resultid="4611" />
                    <RANKING order="30" place="30" resultid="2829" />
                    <RANKING order="31" place="31" resultid="3308" />
                    <RANKING order="32" place="32" resultid="2684" />
                    <RANKING order="33" place="33" resultid="2966" />
                    <RANKING order="34" place="34" resultid="3667" />
                    <RANKING order="35" place="35" resultid="3867" />
                    <RANKING order="36" place="36" resultid="3888" />
                    <RANKING order="37" place="37" resultid="2676" />
                    <RANKING order="38" place="38" resultid="3156" />
                    <RANKING order="39" place="39" resultid="2554" />
                    <RANKING order="40" place="40" resultid="2877" />
                    <RANKING order="41" place="41" resultid="3363" />
                    <RANKING order="42" place="42" resultid="4028" />
                    <RANKING order="43" place="43" resultid="2836" />
                    <RANKING order="44" place="44" resultid="2424" />
                    <RANKING order="45" place="45" resultid="4104" />
                    <RANKING order="46" place="46" resultid="3324" />
                    <RANKING order="47" place="47" resultid="3101" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4709" daytime="11:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4710" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4711" daytime="11:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4712" daytime="11:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4713" daytime="11:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4714" daytime="11:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4715" daytime="11:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4716" daytime="11:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5369" gender="M" number="6" order="30" round="SOP" preveventid="1778">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5375" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5377" />
                    <RANKING order="2" place="2" resultid="5376" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5378" agegroupid="5375" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1059" daytime="10:00" gender="F" number="1" order="1" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1060" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3503" />
                    <RANKING order="2" place="2" resultid="3586" />
                    <RANKING order="3" place="3" resultid="2871" />
                    <RANKING order="4" place="4" resultid="2940" />
                    <RANKING order="5" place="5" resultid="3059" />
                    <RANKING order="6" place="6" resultid="3284" />
                    <RANKING order="7" place="7" resultid="4065" />
                    <RANKING order="8" place="8" resultid="3531" />
                    <RANKING order="9" place="9" resultid="3293" />
                    <RANKING order="10" place="10" resultid="3265" />
                    <RANKING order="11" place="11" resultid="2973" />
                    <RANKING order="12" place="12" resultid="3752" />
                    <RANKING order="13" place="13" resultid="2960" />
                    <RANKING order="14" place="14" resultid="3547" />
                    <RANKING order="15" place="15" resultid="3479" />
                    <RANKING order="16" place="16" resultid="4149" />
                    <RANKING order="17" place="17" resultid="2923" />
                    <RANKING order="18" place="17" resultid="3609" />
                    <RANKING order="19" place="19" resultid="3107" />
                    <RANKING order="20" place="20" resultid="3218" />
                    <RANKING order="21" place="21" resultid="2471" />
                    <RANKING order="22" place="22" resultid="3232" />
                    <RANKING order="23" place="23" resultid="3240" />
                    <RANKING order="24" place="24" resultid="3726" />
                    <RANKING order="25" place="25" resultid="4057" />
                    <RANKING order="26" place="26" resultid="4251" />
                    <RANKING order="27" place="27" resultid="3271" />
                    <RANKING order="28" place="28" resultid="3353" />
                    <RANKING order="29" place="29" resultid="2455" />
                    <RANKING order="30" place="29" resultid="3836" />
                    <RANKING order="31" place="31" resultid="2505" />
                    <RANKING order="32" place="32" resultid="3809" />
                    <RANKING order="33" place="33" resultid="3175" />
                    <RANKING order="34" place="34" resultid="3202" />
                    <RANKING order="35" place="35" resultid="2761" />
                    <RANKING order="36" place="36" resultid="3684" />
                    <RANKING order="37" place="37" resultid="3370" />
                    <RANKING order="38" place="38" resultid="3395" />
                    <RANKING order="39" place="39" resultid="2689" />
                    <RANKING order="40" place="39" resultid="3615" />
                    <RANKING order="41" place="41" resultid="2883" />
                    <RANKING order="42" place="42" resultid="3912" />
                    <RANKING order="43" place="43" resultid="4656" />
                    <RANKING order="44" place="44" resultid="2679" />
                    <RANKING order="45" place="45" resultid="4200" />
                    <RANKING order="46" place="46" resultid="3255" />
                    <RANKING order="47" place="47" resultid="4954" />
                    <RANKING order="48" place="48" resultid="3428" />
                    <RANKING order="49" place="49" resultid="2722" />
                    <RANKING order="50" place="50" resultid="4108" />
                    <RANKING order="51" place="51" resultid="3047" />
                    <RANKING order="52" place="52" resultid="2744" />
                    <RANKING order="53" place="53" resultid="2617" />
                    <RANKING order="54" place="54" resultid="3735" />
                    <RANKING order="55" place="55" resultid="3333" />
                    <RANKING order="56" place="56" resultid="2865" />
                    <RANKING order="57" place="57" resultid="3115" />
                    <RANKING order="58" place="58" resultid="4051" />
                    <RANKING order="59" place="59" resultid="2576" />
                    <RANKING order="60" place="59" resultid="3419" />
                    <RANKING order="61" place="61" resultid="2594" />
                    <RANKING order="62" place="62" resultid="4261" />
                    <RANKING order="63" place="63" resultid="2753" />
                    <RANKING order="64" place="64" resultid="4220" />
                    <RANKING order="65" place="65" resultid="2519" />
                    <RANKING order="66" place="66" resultid="2527" />
                    <RANKING order="67" place="66" resultid="3225" />
                    <RANKING order="68" place="68" resultid="3382" />
                    <RANKING order="69" place="69" resultid="3681" />
                    <RANKING order="70" place="70" resultid="2986" />
                    <RANKING order="71" place="71" resultid="3920" />
                    <RANKING order="72" place="72" resultid="2713" />
                    <RANKING order="73" place="73" resultid="4227" />
                    <RANKING order="74" place="74" resultid="3003" />
                    <RANKING order="75" place="75" resultid="4003" />
                    <RANKING order="76" place="76" resultid="4135" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4662" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4663" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4664" daytime="10:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4665" daytime="10:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4666" daytime="10:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4667" daytime="10:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4668" daytime="10:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4669" daytime="10:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4670" daytime="10:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4671" daytime="10:10" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4672" daytime="10:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4673" daytime="10:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4674" daytime="10:15" number="13" order="13" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5443" gender="M" number="14" order="31" round="SOP" preveventid="1834">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5449" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5450" />
                    <RANKING order="2" place="2" resultid="5451" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5452" agegroupid="5449" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1848" daytime="14:25" gender="M" number="16" order="27" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1849" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2968" />
                    <RANKING order="2" place="2" resultid="2607" />
                    <RANKING order="3" place="3" resultid="4236" />
                    <RANKING order="4" place="4" resultid="3623" />
                    <RANKING order="5" place="5" resultid="3476" />
                    <RANKING order="6" place="6" resultid="3130" />
                    <RANKING order="7" place="7" resultid="3526" />
                    <RANKING order="8" place="8" resultid="4184" />
                    <RANKING order="9" place="9" resultid="3054" />
                    <RANKING order="10" place="10" resultid="3190" />
                    <RANKING order="11" place="11" resultid="3984" />
                    <RANKING order="12" place="12" resultid="3443" />
                    <RANKING order="13" place="13" resultid="3935" />
                    <RANKING order="14" place="14" resultid="2416" />
                    <RANKING order="15" place="15" resultid="4119" />
                    <RANKING order="16" place="16" resultid="3714" />
                    <RANKING order="17" place="17" resultid="4176" />
                    <RANKING order="18" place="18" resultid="2781" />
                    <RANKING order="19" place="19" resultid="2706" />
                    <RANKING order="20" place="20" resultid="2556" />
                    <RANKING order="21" place="21" resultid="2843" />
                    <RANKING order="22" place="22" resultid="3777" />
                    <RANKING order="23" place="23" resultid="3168" />
                    <RANKING order="24" place="24" resultid="3890" />
                    <RANKING order="25" place="25" resultid="3762" />
                    <RANKING order="26" place="26" resultid="2538" />
                    <RANKING order="27" place="27" resultid="3289" />
                    <RANKING order="28" place="28" resultid="2732" />
                    <RANKING order="29" place="29" resultid="4030" />
                    <RANKING order="30" place="30" resultid="3904" />
                    <RANKING order="31" place="31" resultid="3972" />
                    <RANKING order="32" place="32" resultid="3309" />
                    <RANKING order="33" place="33" resultid="2647" />
                    <RANKING order="34" place="34" resultid="2654" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4786" daytime="14:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4787" daytime="14:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4788" daytime="14:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4789" daytime="14:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4790" daytime="14:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4791" daytime="14:35" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1771" daytime="11:00" gender="F" number="5" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1772" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3604" />
                    <RANKING order="2" place="2" resultid="3964" />
                    <RANKING order="3" place="3" resultid="3580" />
                    <RANKING order="4" place="4" resultid="2961" />
                    <RANKING order="5" place="5" resultid="4194" />
                    <RANKING order="6" place="6" resultid="2562" />
                    <RANKING order="7" place="7" resultid="3149" />
                    <RANKING order="8" place="8" resultid="3977" />
                    <RANKING order="9" place="9" resultid="3537" />
                    <RANKING order="10" place="10" resultid="3719" />
                    <RANKING order="11" place="11" resultid="3067" />
                    <RANKING order="12" place="12" resultid="4210" />
                    <RANKING order="13" place="13" resultid="4597" />
                    <RANKING order="14" place="14" resultid="3041" />
                    <RANKING order="15" place="15" resultid="4228" />
                    <RANKING order="16" place="16" resultid="3952" />
                    <RANKING order="17" place="17" resultid="3305" />
                    <RANKING order="18" place="18" resultid="4005" />
                    <RANKING order="19" place="19" resultid="3233" />
                    <RANKING order="20" place="-1" resultid="3575" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4705" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4706" daytime="11:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4707" daytime="11:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4708" daytime="11:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1855" daytime="14:40" gender="F" number="17" order="28" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1856" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2994" />
                    <RANKING order="2" place="2" resultid="3593" />
                    <RANKING order="3" place="3" resultid="3928" />
                    <RANKING order="4" place="4" resultid="2873" />
                    <RANKING order="5" place="5" resultid="3533" />
                    <RANKING order="6" place="6" resultid="2974" />
                    <RANKING order="7" place="7" resultid="3286" />
                    <RANKING order="8" place="8" resultid="2671" />
                    <RANKING order="9" place="9" resultid="4168" />
                    <RANKING order="10" place="10" resultid="4153" />
                    <RANKING order="11" place="11" resultid="3355" />
                    <RANKING order="12" place="12" resultid="3016" />
                    <RANKING order="13" place="13" resultid="3803" />
                    <RANKING order="14" place="14" resultid="3727" />
                    <RANKING order="15" place="15" resultid="3272" />
                    <RANKING order="16" place="16" resultid="2457" />
                    <RANKING order="17" place="16" resultid="3258" />
                    <RANKING order="18" place="18" resultid="3144" />
                    <RANKING order="19" place="19" resultid="3024" />
                    <RANKING order="20" place="20" resultid="2487" />
                    <RANKING order="21" place="21" resultid="3947" />
                    <RANKING order="22" place="22" resultid="4059" />
                    <RANKING order="23" place="23" resultid="2796" />
                    <RANKING order="24" place="24" resultid="2596" />
                    <RANKING order="25" place="24" resultid="4252" />
                    <RANKING order="26" place="26" resultid="2578" />
                    <RANKING order="27" place="27" resultid="4110" />
                    <RANKING order="28" place="28" resultid="4652" />
                    <RANKING order="29" place="29" resultid="3372" />
                    <RANKING order="30" place="30" resultid="3431" />
                    <RANKING order="31" place="31" resultid="3243" />
                    <RANKING order="32" place="32" resultid="4196" />
                    <RANKING order="33" place="33" resultid="3438" />
                    <RANKING order="34" place="34" resultid="4081" />
                    <RANKING order="35" place="35" resultid="2543" />
                    <RANKING order="36" place="35" resultid="2680" />
                    <RANKING order="37" place="35" resultid="3221" />
                    <RANKING order="38" place="38" resultid="4580" />
                    <RANKING order="39" place="39" resultid="4046" />
                    <RANKING order="40" place="39" resultid="4658" />
                    <RANKING order="41" place="41" resultid="4076" />
                    <RANKING order="42" place="42" resultid="3721" />
                    <RANKING order="43" place="43" resultid="3682" />
                    <RANKING order="44" place="44" resultid="2935" />
                    <RANKING order="45" place="44" resultid="3954" />
                    <RANKING order="46" place="46" resultid="2619" />
                    <RANKING order="47" place="47" resultid="4956" />
                    <RANKING order="48" place="48" resultid="2697" />
                    <RANKING order="49" place="49" resultid="4007" />
                    <RANKING order="50" place="50" resultid="3185" />
                    <RANKING order="51" place="51" resultid="2867" />
                    <RANKING order="52" place="52" resultid="2769" />
                    <RANKING order="53" place="53" resultid="3845" />
                    <RANKING order="54" place="-1" resultid="3033" />
                    <RANKING order="55" place="-1" resultid="3878" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4793" daytime="14:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4794" daytime="14:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4795" daytime="14:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4796" daytime="14:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4797" daytime="14:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4798" daytime="14:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4799" daytime="14:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4800" daytime="14:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4801" daytime="14:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4961" daytime="14:45" number="10" order="10" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1799" daytime="12:25" gender="F" number="9" order="16" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1800" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3592" />
                    <RANKING order="2" place="2" resultid="3143" />
                    <RANKING order="3" place="3" resultid="3833" />
                    <RANKING order="4" place="4" resultid="2993" />
                    <RANKING order="5" place="5" resultid="2872" />
                    <RANKING order="6" place="6" resultid="3285" />
                    <RANKING order="7" place="7" resultid="3860" />
                    <RANKING order="8" place="8" resultid="3300" />
                    <RANKING order="9" place="9" resultid="4044" />
                    <RANKING order="10" place="10" resultid="4257" />
                    <RANKING order="11" place="11" resultid="2473" />
                    <RANKING order="12" place="12" resultid="3176" />
                    <RANKING order="13" place="13" resultid="2670" />
                    <RANKING order="14" place="14" resultid="3430" />
                    <RANKING order="15" place="15" resultid="4109" />
                    <RANKING order="16" place="16" resultid="4152" />
                    <RANKING order="17" place="17" resultid="2763" />
                    <RANKING order="18" place="18" resultid="3414" />
                    <RANKING order="19" place="19" resultid="2815" />
                    <RANKING order="20" place="20" resultid="2486" />
                    <RANKING order="21" place="21" resultid="3437" />
                    <RANKING order="22" place="22" resultid="2746" />
                    <RANKING order="23" place="23" resultid="3256" />
                    <RANKING order="24" place="24" resultid="2478" />
                    <RANKING order="25" place="25" resultid="2542" />
                    <RANKING order="26" place="26" resultid="3371" />
                    <RANKING order="27" place="27" resultid="2618" />
                    <RANKING order="28" place="28" resultid="3420" />
                    <RANKING order="29" place="29" resultid="3220" />
                    <RANKING order="30" place="30" resultid="2795" />
                    <RANKING order="31" place="31" resultid="4651" />
                    <RANKING order="32" place="32" resultid="3042" />
                    <RANKING order="33" place="33" resultid="3241" />
                    <RANKING order="34" place="34" resultid="4013" />
                    <RANKING order="35" place="35" resultid="2508" />
                    <RANKING order="36" place="36" resultid="3387" />
                    <RANKING order="37" place="37" resultid="2716" />
                    <RANKING order="38" place="38" resultid="2595" />
                    <RANKING order="39" place="39" resultid="4657" />
                    <RANKING order="40" place="40" resultid="2448" />
                    <RANKING order="41" place="41" resultid="2723" />
                    <RANKING order="42" place="42" resultid="3068" />
                    <RANKING order="43" place="43" resultid="3005" />
                    <RANKING order="44" place="44" resultid="3234" />
                    <RANKING order="45" place="45" resultid="3306" />
                    <RANKING order="46" place="46" resultid="2521" />
                    <RANKING order="47" place="47" resultid="2754" />
                    <RANKING order="48" place="48" resultid="2768" />
                    <RANKING order="49" place="49" resultid="2529" />
                    <RANKING order="50" place="50" resultid="3227" />
                    <RANKING order="51" place="51" resultid="3184" />
                    <RANKING order="52" place="-1" resultid="3876" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4728" daytime="12:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4729" daytime="12:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4730" daytime="12:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4731" daytime="12:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4732" daytime="12:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4733" daytime="12:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4734" daytime="12:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4735" daytime="12:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4736" daytime="12:35" number="9" order="9" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1834" daytime="13:55" gender="M" number="14" order="24" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1835" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3038" />
                    <RANKING order="2" place="2" resultid="3598" />
                    <RANKING order="3" place="3" resultid="3195" />
                    <RANKING order="4" place="4" resultid="3989" />
                    <RANKING order="5" place="5" resultid="3564" />
                    <RANKING order="6" place="6" resultid="3676" />
                    <RANKING order="7" place="7" resultid="4224" />
                    <RANKING order="8" place="8" resultid="3698" />
                    <RANKING order="9" place="9" resultid="3983" />
                    <RANKING order="10" place="10" resultid="3692" />
                    <RANKING order="11" place="11" resultid="2799" />
                    <RANKING order="12" place="12" resultid="3510" />
                    <RANKING order="13" place="13" resultid="2441" />
                    <RANKING order="14" place="13" resultid="3277" />
                    <RANKING order="15" place="15" resultid="3137" />
                    <RANKING order="16" place="16" resultid="3467" />
                    <RANKING order="17" place="17" resultid="3499" />
                    <RANKING order="18" place="18" resultid="4215" />
                    <RANKING order="19" place="19" resultid="2451" />
                    <RANKING order="20" place="20" resultid="2854" />
                    <RANKING order="21" place="21" resultid="2819" />
                    <RANKING order="22" place="22" resultid="3662" />
                    <RANKING order="23" place="23" resultid="2998" />
                    <RANKING order="24" place="24" resultid="4139" />
                    <RANKING order="25" place="25" resultid="3348" />
                    <RANKING order="26" place="26" resultid="2892" />
                    <RANKING order="27" place="27" resultid="4183" />
                    <RANKING order="28" place="28" resultid="2685" />
                    <RANKING order="29" place="28" resultid="3873" />
                    <RANKING order="30" place="30" resultid="3082" />
                    <RANKING order="31" place="31" resultid="3365" />
                    <RANKING order="32" place="32" resultid="2633" />
                    <RANKING order="33" place="32" resultid="3668" />
                    <RANKING order="34" place="34" resultid="2626" />
                    <RANKING order="35" place="35" resultid="2848" />
                    <RANKING order="36" place="35" resultid="2980" />
                    <RANKING order="37" place="37" resultid="3102" />
                    <RANKING order="38" place="38" resultid="2954" />
                    <RANKING order="39" place="39" resultid="3732" />
                    <RANKING order="40" place="40" resultid="3658" />
                    <RANKING order="41" place="41" resultid="3853" />
                    <RANKING order="42" place="42" resultid="2426" />
                    <RANKING order="43" place="42" resultid="4021" />
                    <RANKING order="44" place="44" resultid="3903" />
                    <RANKING order="45" place="45" resultid="3401" />
                    <RANKING order="46" place="46" resultid="2842" />
                    <RANKING order="47" place="47" resultid="3490" />
                    <RANKING order="48" place="48" resultid="3868" />
                    <RANKING order="49" place="49" resultid="2823" />
                    <RANKING order="50" place="50" resultid="2898" />
                    <RANKING order="51" place="51" resultid="3450" />
                    <RANKING order="52" place="52" resultid="2667" />
                    <RANKING order="53" place="52" resultid="3748" />
                    <RANKING order="54" place="54" resultid="3883" />
                    <RANKING order="55" place="55" resultid="3743" />
                    <RANKING order="56" place="56" resultid="4587" />
                    <RANKING order="57" place="57" resultid="3456" />
                    <RANKING order="58" place="58" resultid="3521" />
                    <RANKING order="59" place="59" resultid="2409" />
                    <RANKING order="60" place="60" resultid="4642" />
                    <RANKING order="61" place="61" resultid="2878" />
                    <RANKING order="62" place="62" resultid="2807" />
                    <RANKING order="63" place="63" resultid="3361" />
                    <RANKING order="64" place="64" resultid="4570" />
                    <RANKING order="65" place="65" resultid="2537" />
                    <RANKING order="66" place="66" resultid="4638" />
                    <RANKING order="67" place="67" resultid="2493" />
                    <RANKING order="68" place="68" resultid="2661" />
                    <RANKING order="69" place="69" resultid="2404" />
                    <RANKING order="70" place="70" resultid="2739" />
                    <RANKING order="71" place="71" resultid="2584" />
                    <RANKING order="72" place="-1" resultid="2641" />
                    <RANKING order="73" place="-1" resultid="3158" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4765" daytime="13:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4766" daytime="13:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4767" daytime="13:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4768" daytime="13:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4769" daytime="13:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4770" daytime="13:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4771" daytime="13:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4772" daytime="14:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4773" daytime="14:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4774" daytime="14:00" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4775" daytime="14:00" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4776" daytime="14:00" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4777" daytime="14:00" number="13" order="13" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-11-05" daytime="16:45" endtime="19:39" number="2">
          <EVENTS>
            <EVENT eventid="1919" gender="F" number="9" order="25" round="FIN" preveventid="1799">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1920" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5392" />
                    <RANKING order="2" place="2" resultid="5395" />
                    <RANKING order="3" place="3" resultid="5393" />
                    <RANKING order="4" place="4" resultid="5394" />
                    <RANKING order="5" place="5" resultid="5396" />
                    <RANKING order="6" place="6" resultid="5397" />
                    <RANKING order="7" place="7" resultid="5399" />
                    <RANKING order="8" place="8" resultid="5398" />
                    <RANKING order="9" place="9" resultid="5401" />
                    <RANKING order="10" place="10" resultid="5400" />
                    <RANKING order="11" place="11" resultid="5403" />
                    <RANKING order="12" place="12" resultid="5402" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5404" agegroupid="1920" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4737" agegroupid="1920" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1898" gender="M" number="6" order="18" round="FIN" preveventid="1778">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1899" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5453" />
                    <RANKING order="2" place="2" resultid="5454" />
                    <RANKING order="3" place="3" resultid="5457" />
                    <RANKING order="4" place="4" resultid="5458" />
                    <RANKING order="5" place="5" resultid="5455" />
                    <RANKING order="6" place="6" resultid="5456" />
                    <RANKING order="7" place="7" resultid="5461" />
                    <RANKING order="8" place="8" resultid="5460" />
                    <RANKING order="9" place="9" resultid="5462" />
                    <RANKING order="10" place="10" resultid="5463" />
                    <RANKING order="11" place="11" resultid="5459" />
                    <RANKING order="12" place="12" resultid="5464" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5465" agegroupid="1899" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4717" agegroupid="1899" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1905" gender="F" number="18" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1906" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3588" />
                    <RANKING order="2" place="2" resultid="3549" />
                    <RANKING order="3" place="3" resultid="3539" />
                    <RANKING order="4" place="4" resultid="3611" />
                    <RANKING order="5" place="5" resultid="3582" />
                    <RANKING order="6" place="6" resultid="3178" />
                    <RANKING order="7" place="7" resultid="3755" />
                    <RANKING order="8" place="8" resultid="3838" />
                    <RANKING order="9" place="9" resultid="4230" />
                    <RANKING order="10" place="10" resultid="3049" />
                    <RANKING order="11" place="11" resultid="3117" />
                    <RANKING order="12" place="12" resultid="3722" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4803" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4804" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1863" gender="F" number="1" order="3" round="FIN" preveventid="1059">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1864" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="5318" />
                    <RANKING order="2" place="-1" resultid="5319" />
                    <RANKING order="3" place="-1" resultid="5320" />
                    <RANKING order="4" place="-1" resultid="5323" />
                    <RANKING order="5" place="-1" resultid="5321" />
                    <RANKING order="6" place="-1" resultid="5322" />
                    <RANKING order="7" place="-1" resultid="5325" />
                    <RANKING order="8" place="-1" resultid="5324" />
                    <RANKING order="9" place="-1" resultid="5327" />
                    <RANKING order="10" place="-1" resultid="5326" />
                    <RANKING order="11" place="-1" resultid="5329" />
                    <RANKING order="12" place="-1" resultid="5328" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5317" agegroupid="1864" final="B" number="1" order="1" status="INOFFICIAL" />
                <HEAT heatid="4675" agegroupid="1864" final="A" number="2" order="2" status="INOFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1926" gender="M" number="12" order="27" round="FIN" preveventid="1820">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1927" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5430" />
                    <RANKING order="2" place="2" resultid="5432" />
                    <RANKING order="3" place="3" resultid="5433" />
                    <RANKING order="4" place="4" resultid="5431" />
                    <RANKING order="5" place="5" resultid="5434" />
                    <RANKING order="6" place="6" resultid="5435" />
                    <RANKING order="7" place="7" resultid="5438" />
                    <RANKING order="8" place="8" resultid="5436" />
                    <RANKING order="9" place="9" resultid="5439" />
                    <RANKING order="10" place="10" resultid="5441" />
                    <RANKING order="11" place="11" resultid="5440" />
                    <RANKING order="12" place="12" resultid="5437" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5442" agegroupid="1927" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4757" agegroupid="1927" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1954" gender="F" number="15" order="33" round="FIN" preveventid="1841">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1955" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5479" />
                    <RANKING order="2" place="2" resultid="5480" />
                    <RANKING order="3" place="3" resultid="5481" />
                    <RANKING order="4" place="4" resultid="5482" />
                    <RANKING order="5" place="5" resultid="5484" />
                    <RANKING order="6" place="6" resultid="5483" />
                    <RANKING order="7" place="7" resultid="5487" />
                    <RANKING order="8" place="8" resultid="5486" />
                    <RANKING order="9" place="9" resultid="5489" />
                    <RANKING order="10" place="10" resultid="5488" />
                    <RANKING order="11" place="11" resultid="5485" />
                    <RANKING order="12" place="12" resultid="5490" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5491" agegroupid="1955" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4785" agegroupid="1955" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1884" gender="M" number="4" order="13" round="FIN" preveventid="1763">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1885" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5356" />
                    <RANKING order="2" place="2" resultid="5357" />
                    <RANKING order="3" place="3" resultid="5358" />
                    <RANKING order="4" place="4" resultid="5360" />
                    <RANKING order="5" place="5" resultid="5359" />
                    <RANKING order="6" place="6" resultid="5361" />
                    <RANKING order="7" place="7" resultid="5363" />
                    <RANKING order="8" place="8" resultid="5362" />
                    <RANKING order="9" place="9" resultid="5364" />
                    <RANKING order="10" place="10" resultid="5366" />
                    <RANKING order="11" place="11" resultid="5365" />
                    <RANKING order="12" place="-1" resultid="5367" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5368" agegroupid="1885" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4704" agegroupid="1885" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2062" gender="F" number="20" order="41" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="2000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2063" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3638" />
                    <RANKING order="2" place="2" resultid="3199" />
                    <RANKING order="3" place="3" resultid="4085" />
                    <RANKING order="4" place="4" resultid="2904" />
                    <RANKING order="5" place="5" resultid="3327" />
                    <RANKING order="6" place="6" resultid="3783" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4807" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1870" gender="M" number="2" order="6" round="FIN" preveventid="1749">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="5342" agegroupid="1871" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4686" agegroupid="1871" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1891" gender="F" number="7" order="15" round="FIN" preveventid="1785">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1892" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5382" />
                    <RANKING order="2" place="2" resultid="5379" />
                    <RANKING order="3" place="3" resultid="5380" />
                    <RANKING order="4" place="4" resultid="5381" />
                    <RANKING order="5" place="5" resultid="5383" />
                    <RANKING order="6" place="6" resultid="5384" />
                    <RANKING order="7" place="7" resultid="5385" />
                    <RANKING order="8" place="8" resultid="5387" />
                    <RANKING order="9" place="9" resultid="5386" />
                    <RANKING order="10" place="10" resultid="5390" />
                    <RANKING order="11" place="11" resultid="5388" />
                    <RANKING order="12" place="12" resultid="5389" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5391" agegroupid="1892" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4725" agegroupid="1892" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1912" gender="M" number="10" order="23" round="FIN" preveventid="1806">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1913" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5405" />
                    <RANKING order="2" place="2" resultid="5406" />
                    <RANKING order="3" place="3" resultid="5408" />
                    <RANKING order="4" place="4" resultid="5407" />
                    <RANKING order="5" place="5" resultid="5410" />
                    <RANKING order="6" place="6" resultid="5409" />
                    <RANKING order="7" place="7" resultid="5411" />
                    <RANKING order="8" place="8" resultid="5413" />
                    <RANKING order="9" place="9" resultid="5412" />
                    <RANKING order="10" place="10" resultid="5414" />
                    <RANKING order="11" place="11" resultid="5415" />
                    <RANKING order="12" place="12" resultid="5416" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5417" agegroupid="1913" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4744" agegroupid="1913" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1947" gender="M" number="14" order="31" round="FIN" preveventid="1834">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1948" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5466" />
                    <RANKING order="2" place="2" resultid="5467" />
                    <RANKING order="3" place="3" resultid="5468" />
                    <RANKING order="4" place="4" resultid="5469" />
                    <RANKING order="5" place="5" resultid="5470" />
                    <RANKING order="6" place="6" resultid="5471" />
                    <RANKING order="7" place="7" resultid="5472" />
                    <RANKING order="8" place="8" resultid="5475" />
                    <RANKING order="9" place="9" resultid="5477" />
                    <RANKING order="10" place="10" resultid="5474" />
                    <RANKING order="11" place="11" resultid="5476" />
                    <RANKING order="12" place="12" resultid="5473" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5478" agegroupid="1948" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4778" agegroupid="1948" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1961" gender="M" number="16" order="35" round="FIN" preveventid="1848">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1962" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5492" />
                    <RANKING order="2" place="2" resultid="5493" />
                    <RANKING order="3" place="3" resultid="5494" />
                    <RANKING order="4" place="4" resultid="5495" />
                    <RANKING order="5" place="5" resultid="5497" />
                    <RANKING order="6" place="6" resultid="5496" />
                    <RANKING order="7" place="7" resultid="5499" />
                    <RANKING order="8" place="8" resultid="5498" />
                    <RANKING order="9" place="9" resultid="5500" />
                    <RANKING order="10" place="10" resultid="5503" />
                    <RANKING order="11" place="11" resultid="5502" />
                    <RANKING order="12" place="12" resultid="5501" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5504" agegroupid="1962" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4792" agegroupid="1962" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1877" gender="F" number="3" order="10" round="FIN" preveventid="1756">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1878" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5343" />
                    <RANKING order="2" place="2" resultid="5348" />
                    <RANKING order="3" place="3" resultid="5345" />
                    <RANKING order="4" place="4" resultid="5346" />
                    <RANKING order="5" place="5" resultid="5344" />
                    <RANKING order="6" place="6" resultid="5347" />
                    <RANKING order="7" place="7" resultid="5352" />
                    <RANKING order="8" place="8" resultid="5353" />
                    <RANKING order="9" place="9" resultid="5351" />
                    <RANKING order="10" place="10" resultid="5349" />
                    <RANKING order="11" place="11" resultid="5350" />
                    <RANKING order="12" place="12" resultid="5354" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5355" agegroupid="1878" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4695" agegroupid="1878" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2048" gender="M" number="19" order="40" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="2000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2396" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3197" />
                    <RANKING order="2" place="2" resultid="3636" />
                    <RANKING order="3" place="3" resultid="4083" />
                    <RANKING order="4" place="4" resultid="4240" />
                    <RANKING order="5" place="5" resultid="4158" />
                    <RANKING order="6" place="6" resultid="3702" />
                    <RANKING order="7" place="7" resultid="3492" />
                    <RANKING order="8" place="8" resultid="4626" />
                    <RANKING order="9" place="9" resultid="3781" />
                    <RANKING order="10" place="-1" resultid="2902" />
                    <RANKING order="11" place="-1" resultid="3704" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4805" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4806" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1933" gender="F" number="11" order="29" round="FIN" preveventid="1813">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1934" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5418" />
                    <RANKING order="2" place="2" resultid="5419" />
                    <RANKING order="3" place="3" resultid="5421" />
                    <RANKING order="4" place="4" resultid="5423" />
                    <RANKING order="5" place="5" resultid="5422" />
                    <RANKING order="6" place="6" resultid="5420" />
                    <RANKING order="7" place="7" resultid="5426" />
                    <RANKING order="8" place="8" resultid="5427" />
                    <RANKING order="9" place="9" resultid="5425" />
                    <RANKING order="10" place="10" resultid="5424" />
                    <RANKING order="11" place="11" resultid="5428" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5429" agegroupid="1934" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4748" agegroupid="1934" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1940" gender="F" number="17" order="37" round="FIN" preveventid="1855">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1941" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5505" />
                    <RANKING order="2" place="2" resultid="5506" />
                    <RANKING order="3" place="3" resultid="5508" />
                    <RANKING order="4" place="4" resultid="5507" />
                    <RANKING order="5" place="5" resultid="5509" />
                    <RANKING order="6" place="6" resultid="5510" />
                    <RANKING order="7" place="7" resultid="5513" />
                    <RANKING order="8" place="8" resultid="5511" />
                    <RANKING order="9" place="9" resultid="5514" />
                    <RANKING order="10" place="10" resultid="5515" />
                    <RANKING order="11" place="11" resultid="5512" />
                    <RANKING order="12" place="12" resultid="5516" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5517" agegroupid="1941" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4802" agegroupid="1941" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-11-06" daytime="09:30" number="3" officialmeeting="09:00" teamleadermeeting="09:00" warmupfrom="07:45" warmupuntil="09:15">
          <EVENTS>
            <EVENT eventid="1999" daytime="10:35" gender="M" number="25" order="32" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4859" daytime="10:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4860" daytime="10:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4861" daytime="10:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4862" daytime="10:50" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1971" daytime="09:30" gender="M" number="21" order="23" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4813" daytime="09:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4814" daytime="09:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4815" daytime="09:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4816" daytime="09:35" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4817" daytime="09:35" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4818" daytime="09:35" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4819" daytime="09:35" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4820" daytime="09:40" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4821" daytime="09:40" number="9" order="9" status="SEEDED" />
                <HEAT heatid="4822" daytime="09:40" number="10" order="10" status="SEEDED" />
                <HEAT heatid="4823" daytime="09:40" number="11" order="11" status="SEEDED" />
                <HEAT heatid="4824" daytime="09:45" number="12" order="12" status="SEEDED" />
                <HEAT heatid="4825" daytime="09:45" number="13" order="13" status="SEEDED" />
                <HEAT heatid="4826" daytime="09:45" number="14" order="14" status="SEEDED" />
                <HEAT heatid="4827" daytime="09:45" number="15" order="15" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2096" daytime="13:30" gender="F" number="36" order="49" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4932" daytime="13:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4933" daytime="13:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4934" daytime="13:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4935" daytime="13:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4936" daytime="13:40" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4937" daytime="13:45" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1985" daytime="10:15" gender="M" number="23" order="28" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4840" daytime="10:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4841" daytime="10:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4842" daytime="10:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4843" daytime="10:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4844" daytime="10:20" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4845" daytime="10:20" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4846" daytime="10:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4847" daytime="10:20" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4848" daytime="10:20" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2027" daytime="11:35" gender="M" number="29" order="39" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4877" daytime="11:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4878" daytime="11:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4879" daytime="11:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4880" daytime="11:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4881" daytime="11:40" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2013" daytime="11:05" gender="M" number="27" order="36" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2014" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4237" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4869" daytime="11:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4870" daytime="11:10" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4871" daytime="11:10" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4872" daytime="11:10" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4873" daytime="11:10" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1978" daytime="09:50" gender="F" number="22" order="26" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4829" daytime="09:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4830" daytime="09:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4831" daytime="09:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4832" daytime="09:55" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4833" daytime="10:00" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4834" daytime="10:00" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4835" daytime="10:05" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4836" daytime="10:05" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4837" daytime="10:10" number="9" order="9" status="SEEDED" />
                <HEAT heatid="4838" daytime="10:10" number="10" order="10" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1992" daytime="10:20" gender="F" number="24" order="30" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4850" daytime="10:20" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4851" daytime="10:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4852" daytime="10:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4853" daytime="10:25" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4854" daytime="10:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4855" daytime="10:30" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4856" daytime="10:30" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4857" daytime="10:35" number="8" order="8" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2055" daytime="12:00" gender="F" number="32" order="43" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4896" daytime="12:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4897" daytime="12:05" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4898" daytime="12:10" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4899" daytime="12:10" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4900" daytime="12:15" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4901" daytime="12:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4902" daytime="12:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4903" daytime="12:20" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4904" daytime="12:25" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2075" daytime="12:30" gender="M" number="33" order="44" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4906" daytime="12:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4907" daytime="12:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4908" daytime="12:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4909" daytime="12:45" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4910" daytime="12:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4911" daytime="12:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4912" daytime="12:55" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2034" daytime="11:45" gender="F" number="30" order="41" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4883" daytime="11:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4884" daytime="11:45" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4885" daytime="11:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4886" daytime="11:45" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4887" daytime="11:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4888" daytime="11:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4889" daytime="11:50" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2103" daytime="13:45" gender="M" number="37" order="50" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2104" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4239" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4939" daytime="13:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4940" daytime="13:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4941" daytime="13:50" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4942" daytime="13:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4943" daytime="13:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4944" daytime="13:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4945" daytime="13:50" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4946" daytime="13:50" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4947" daytime="13:55" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2006" daytime="10:55" gender="F" number="26" order="34" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4863" daytime="10:55" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4864" daytime="11:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4865" daytime="11:00" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4866" daytime="11:00" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4867" daytime="11:05" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2041" daytime="11:50" gender="M" number="31" order="42" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2042" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4238" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4891" daytime="11:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4892" daytime="11:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4893" daytime="11:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4894" daytime="12:00" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2082" daytime="13:00" gender="F" number="34" order="46" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4913" daytime="13:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4914" daytime="13:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4915" daytime="13:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4916" daytime="13:05" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4917" daytime="13:05" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4918" daytime="13:05" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4919" daytime="13:05" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4920" daytime="13:05" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4921" daytime="13:05" number="9" order="9" status="SEEDED" />
                <HEAT heatid="4922" daytime="13:10" number="10" order="10" status="SEEDED" />
                <HEAT heatid="4923" daytime="13:10" number="11" order="11" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2089" daytime="13:10" gender="M" number="35" order="48" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4925" daytime="13:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4926" daytime="13:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4927" daytime="13:20" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4928" daytime="13:20" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4929" daytime="13:25" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4930" daytime="13:25" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2020" daytime="11:15" gender="F" number="28" order="37" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4875" daytime="11:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4876" daytime="11:25" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-11-06" daytime="16:00" number="4">
          <EVENTS>
            <EVENT eventid="2154" gender="F" number="26" order="52" round="FIN" preveventid="2006">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="4868" agegroupid="2155" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2210" gender="M" number="35" order="70" round="FIN" preveventid="2089">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="4931" agegroupid="2211" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2168" gender="M" number="38" order="55" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4808" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4809" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2189" gender="M" number="31" order="66" round="FIN" preveventid="2041">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="4895" agegroupid="2190" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2182" gender="F" number="30" order="57" round="FIN" preveventid="2034">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="4890" agegroupid="2183" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2126" gender="M" number="21" order="41" round="FIN" preveventid="1971">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="4828" agegroupid="2127" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2147" gender="F" number="24" order="48" round="FIN" preveventid="1992">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="4858" agegroupid="2148" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2224" gender="F" number="39" order="77" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE value="2000" />
              <HEATS>
                <HEAT heatid="4810" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2133" gender="F" number="22" order="43" round="FIN" preveventid="1978">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="4839" agegroupid="2134" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2112" gender="M" number="37" order="74" round="FIN" preveventid="2103">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="4948" agegroupid="2113" final="A" number="1" order="1" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2175" gender="M" number="29" order="60" round="FIN" preveventid="2027">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="4882" agegroupid="2176" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2232" gender="M" number="40" order="78" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE value="2000" />
              <HEATS>
                <HEAT heatid="4811" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4812" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2140" gender="M" number="23" order="46" round="FIN" preveventid="1985">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="4849" agegroupid="2141" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2203" gender="F" number="34" order="68" round="FIN" preveventid="2082">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="4924" agegroupid="2204" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2196" gender="F" number="32" order="64" round="FIN" preveventid="2055">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="4905" agegroupid="2197" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2217" gender="F" number="36" order="72" round="FIN" preveventid="2096">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="4938" agegroupid="2218" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2161" gender="M" number="27" order="50" round="FIN" preveventid="2013">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="4874" agegroupid="2162" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="4167" nation="GER" region="02" clubid="2398" name="1.SC Schweinfurt">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Daniel" gender="M" lastname="Heidbeck" nation="GER" license="379928" athleteid="2399">
              <RESULTS>
                <RESULT eventid="1763" points="473" swimtime="00:01:11.34" resultid="2400" heatid="4696" lane="4" entrytime="00:01:14.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:34.57" eventid="1985" heatid="4841" lane="1" />
                <ENTRY entrytime="00:02:41.81" eventid="2089" heatid="4925" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Simon" gender="M" lastname="Vollert" nation="GER" license="331888" athleteid="2403">
              <RESULTS>
                <RESULT eventid="1834" points="419" swimtime="00:00:27.06" resultid="2404" heatid="4765" lane="3" entrytime="00:00:27.34" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:34.74" eventid="1985" heatid="4840" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4175" nation="GER" region="02" clubid="2525" name="ASV 1860 Neumarkt">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Anika" gender="F" lastname="Jacksteit" nation="GER" license="266125" athleteid="2526">
              <RESULTS>
                <RESULT eventid="1059" points="484" swimtime="00:01:04.80" resultid="2527" heatid="4665" lane="4" entrytime="00:01:03.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="400" swimtime="00:01:14.64" resultid="2528" heatid="4718" lane="4" entrytime="00:01:13.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="409" swimtime="00:01:16.31" resultid="2529" heatid="4730" lane="5" entrytime="00:01:13.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:33.63" eventid="2034" heatid="4885" lane="1" />
                <ENTRY entrytime="00:00:29.02" eventid="2082" heatid="4916" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4168" nation="GER" region="02" clubid="2759" name="ASV Cham">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Lena" gender="F" lastname="Braun" nation="GER" license="294440" athleteid="2760">
              <RESULTS>
                <RESULT eventid="1059" points="546" swimtime="00:01:02.28" resultid="2761" heatid="4670" lane="1" entrytime="00:01:01.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="509" swimtime="00:00:36.05" resultid="2762" heatid="4694" lane="6" entrytime="00:00:34.84" />
                <RESULT eventid="1799" points="507" swimtime="00:01:11.03" resultid="2763" heatid="4732" lane="5" entrytime="00:01:12.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:18.92" eventid="1992" heatid="4852" lane="3" />
                <ENTRY entrytime="00:00:27.35" eventid="2082" heatid="4921" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Alexandra" gender="F" lastname="Wagner" nation="GER" license="320557" athleteid="2766">
              <RESULTS>
                <RESULT eventid="1756" points="441" swimtime="00:00:37.82" resultid="2767" heatid="4688" lane="3" entrytime="00:00:37.10" />
                <RESULT eventid="1799" points="410" swimtime="00:01:16.27" resultid="2768" heatid="4730" lane="6" entrytime="00:01:14.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="403" swimtime="00:00:32.98" resultid="2769" heatid="4793" lane="4" entrytime="00:00:32.15" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.53" eventid="2082" heatid="4915" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4169" nation="GER" region="02" clubid="4644" name="ATS Kulmbach">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Franz" gender="M" lastname="Prell" nation="GER" license="297312" athleteid="4645">
              <RESULTS>
                <RESULT eventid="1749" points="431" swimtime="00:02:11.49" resultid="4646" heatid="4677" lane="1" entrytime="00:02:09.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="100" swimtime="00:01:02.46" />
                    <SPLIT distance="150" swimtime="00:01:36.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:40.20" eventid="2075" heatid="4906" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4224" nation="GER" region="02" clubid="3447" name="Delphin 77 Herzogenaurach">
          <ATHLETES>
            <ATHLETE birthdate="1992-01-01" firstname="Christian" gender="M" lastname="Ziebuhr" nation="GER" license="139641" athleteid="3448">
              <RESULTS>
                <RESULT eventid="1763" points="490" swimtime="00:01:10.49" resultid="3449" heatid="4700" lane="1" entrytime="00:01:09.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="461" swimtime="00:00:26.22" resultid="3450" heatid="4771" lane="5" entrytime="00:00:25.65" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.35" eventid="1985" heatid="4845" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4233" nation="GER" region="02" clubid="3238" name="DJK Sportbund München">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Stefanie" gender="F" lastname="Ohneiser" nation="GER" license="316235" athleteid="3239">
              <RESULTS>
                <RESULT eventid="1059" points="562" swimtime="00:01:01.67" resultid="3240" heatid="4663" lane="4" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="466" swimtime="00:01:13.05" resultid="3241" heatid="4728" lane="3" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="479" swimtime="00:04:59.57" resultid="3242" heatid="4758" lane="2" entrytime="00:04:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:11.83" />
                    <SPLIT distance="150" swimtime="00:01:50.08" />
                    <SPLIT distance="200" swimtime="00:02:28.23" />
                    <SPLIT distance="250" swimtime="00:03:05.96" />
                    <SPLIT distance="300" swimtime="00:03:44.07" />
                    <SPLIT distance="350" swimtime="00:04:22.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="481" swimtime="00:00:31.10" resultid="3243" heatid="4797" lane="4" entrytime="00:00:31.00" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:18.50" eventid="1978" heatid="4831" lane="4" />
                <ENTRY entrytime="00:02:38.50" eventid="2055" heatid="4898" lane="6" />
                <ENTRY entrytime="00:00:29.50" eventid="2082" heatid="4915" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4300" nation="GER" region="02" clubid="2665" name="SB Bayern 07">
          <ATHLETES>
            <ATHLETE birthdate="1995-01-01" firstname="Tim" gender="M" lastname="Grasser" nation="GER" license="150609" athleteid="2666">
              <RESULTS>
                <RESULT eventid="1834" points="459" swimtime="00:00:26.26" resultid="2667" heatid="4770" lane="4" entrytime="00:00:25.90" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.19" eventid="1971" heatid="4821" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Teresa" gender="F" lastname="Kraus" nation="GER" license="183593" athleteid="2669">
              <RESULTS>
                <RESULT eventid="1799" points="520" swimtime="00:01:10.47" resultid="2670" heatid="4732" lane="4" entrytime="00:01:12.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="569" swimtime="00:00:29.42" resultid="2671" heatid="4961" lane="1" entrytime="00:00:29.68" />
                <RESULT eventid="1919" points="494" swimtime="00:01:11.65" resultid="5403" heatid="5404" lane="6" entrytime="00:01:10.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="571" swimtime="00:00:29.37" resultid="5511" heatid="5517" lane="3" entrytime="00:00:29.42" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:08.50" eventid="2006" heatid="4864" lane="3" />
                <ENTRY entrytime="00:00:29.00" eventid="2082" heatid="4917" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4290" nation="GER" region="02" clubid="2598" name="SC 53 Landshut">
          <ATHLETES>
            <ATHLETE birthdate="1993-01-01" firstname="Verena" gender="F" lastname="Dormehl" nation="GER" license="154254" athleteid="2599">
              <RESULTS>
                <RESULT eventid="1756" points="527" swimtime="00:00:35.65" resultid="2600" heatid="4691" lane="4" entrytime="00:00:35.45" />
                <RESULT eventid="1841" points="514" swimtime="00:02:47.96" resultid="2601" heatid="4781" lane="2" entrytime="00:02:49.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:20.81" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:16.30" eventid="1992" heatid="4856" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Ludwig" gender="M" lastname="Freutsmiedl" nation="GER" license="263873" athleteid="2603">
              <RESULTS>
                <RESULT eventid="1749" points="583" swimtime="00:01:58.95" resultid="2604" heatid="4680" lane="3" entrytime="00:02:02.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="100" swimtime="00:00:57.63" />
                    <SPLIT distance="150" swimtime="00:01:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="504" swimtime="00:00:27.91" resultid="2605" heatid="4743" lane="1" entrytime="00:00:28.65" />
                <RESULT eventid="1820" points="564" swimtime="00:02:12.66" resultid="2606" heatid="4753" lane="5" entrytime="00:02:15.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="100" swimtime="00:01:01.93" />
                    <SPLIT distance="150" swimtime="00:01:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="551" swimtime="00:02:08.84" resultid="2607" heatid="4791" lane="2" entrytime="00:02:11.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:03.23" />
                    <SPLIT distance="150" swimtime="00:01:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1912" points="497" swimtime="00:00:28.05" resultid="5414" heatid="5417" lane="5" entrytime="00:00:27.91" />
                <RESULT eventid="1961" points="564" swimtime="00:02:07.80" resultid="5493" heatid="4792" lane="4" entrytime="00:02:08.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                    <SPLIT distance="150" swimtime="00:01:35.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.44" eventid="1971" heatid="4820" lane="5" />
                <ENTRY entrytime="00:01:01.41" eventid="2013" heatid="4872" lane="5" />
                <ENTRY entrytime="00:04:19.25" eventid="2075" heatid="4910" lane="6" />
                <ENTRY entrytime="00:00:28.63" eventid="2103" heatid="4940" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lena" gender="F" lastname="Köhnke" nation="GER" license="284272" athleteid="2612">
              <RESULTS>
                <RESULT eventid="1756" points="526" swimtime="00:00:35.67" resultid="2613" heatid="4689" lane="5" entrytime="00:00:36.85" />
                <RESULT eventid="1841" points="491" swimtime="00:02:50.55" resultid="2614" heatid="4780" lane="4" entrytime="00:02:53.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:23.38" />
                    <SPLIT distance="150" swimtime="00:02:07.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:19.46" eventid="1992" heatid="4852" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Jana" gender="F" lastname="Lakner" nation="GER" license="281157" athleteid="2616">
              <RESULTS>
                <RESULT eventid="1059" points="516" swimtime="00:01:03.44" resultid="2617" heatid="4666" lane="5" entrytime="00:01:03.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="484" swimtime="00:01:12.17" resultid="2618" heatid="4731" lane="6" entrytime="00:01:12.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="445" swimtime="00:00:31.93" resultid="2619" heatid="4795" lane="6" entrytime="00:00:31.85" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:33.67" eventid="2034" heatid="4885" lane="6" />
                <ENTRY entrytime="00:00:28.45" eventid="2082" heatid="4919" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lukas" gender="M" lastname="Mirsch" nation="GER" license="237415" athleteid="2622">
              <RESULTS>
                <RESULT eventid="1749" points="629" swimtime="00:01:55.93" resultid="2623" heatid="4683" lane="1" entrytime="00:01:56.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="100" swimtime="00:00:57.10" />
                    <SPLIT distance="150" swimtime="00:01:27.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="590" swimtime="00:00:57.73" resultid="2624" heatid="4716" lane="4" entrytime="00:00:57.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="520" swimtime="00:00:27.62" resultid="2625" heatid="4743" lane="4" entrytime="00:00:27.25" />
                <RESULT eventid="1834" points="512" swimtime="00:00:25.32" resultid="2626" heatid="4774" lane="3" entrytime="00:00:24.65" />
                <RESULT eventid="1912" points="476" swimtime="00:00:28.44" resultid="5409" heatid="4744" lane="1" entrytime="00:00:27.62" />
                <RESULT eventid="1898" points="584" swimtime="00:00:57.93" resultid="5455" heatid="4717" lane="2" entrytime="00:00:57.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.82" eventid="1971" heatid="4824" lane="3" />
                <ENTRY entrytime="00:02:06.87" eventid="2041" heatid="4894" lane="4" />
                <ENTRY entrytime="00:00:26.28" eventid="2103" heatid="4946" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Toni" gender="M" lastname="Schmid" nation="GER" license="227470" athleteid="2630">
              <RESULTS>
                <RESULT eventid="1763" points="626" swimtime="00:01:05.00" resultid="2631" heatid="4703" lane="5" entrytime="00:01:04.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="440" swimtime="00:00:29.21" resultid="2632" heatid="4740" lane="5" entrytime="00:00:29.57" />
                <RESULT eventid="1834" points="514" swimtime="00:00:25.28" resultid="2633" heatid="4772" lane="5" entrytime="00:00:25.37" />
                <RESULT eventid="1884" points="608" swimtime="00:01:05.63" resultid="5365" heatid="5368" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.07" eventid="1985" heatid="4848" lane="4" />
                <ENTRY entrytime="00:01:00.70" eventid="2027" heatid="4880" lane="2" />
                <ENTRY entrytime="00:00:27.18" eventid="2103" heatid="4944" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Daniel" gender="M" lastname="Siminenko" nation="GER" license="300185" athleteid="2637">
              <RESULTS>
                <RESULT eventid="1749" status="DNS" swimtime="00:00:00.00" resultid="2638" heatid="4676" lane="2" entrytime="00:02:11.30" />
                <RESULT eventid="1763" status="DNS" swimtime="00:00:00.00" resultid="2639" heatid="4697" lane="6" entrytime="00:01:13.58" />
                <RESULT eventid="1820" status="DNS" swimtime="00:00:00.00" resultid="2640" heatid="4750" lane="5" entrytime="00:02:25.22" />
                <RESULT eventid="1834" status="DNS" swimtime="00:00:00.00" resultid="2641" heatid="4766" lane="3" entrytime="00:00:27.28" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:34.03" eventid="1985" heatid="4841" lane="2" />
                <ENTRY entrytime="00:02:39.38" eventid="2089" heatid="4925" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Tobias" gender="M" lastname="Ulbrich" nation="GER" license="247315" athleteid="2644">
              <RESULTS>
                <RESULT eventid="1749" points="460" swimtime="00:02:08.72" resultid="2645" heatid="4677" lane="3" entrytime="00:02:08.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="100" swimtime="00:01:01.50" />
                    <SPLIT distance="150" swimtime="00:01:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="417" swimtime="00:02:26.67" resultid="2646" heatid="4750" lane="1" entrytime="00:02:25.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="150" swimtime="00:01:53.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="390" swimtime="00:02:24.52" resultid="2647" heatid="4786" lane="5" entrytime="00:02:25.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:47.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:05:08.07" eventid="1999" heatid="4859" lane="2" />
                <ENTRY entrytime="00:04:32.53" eventid="2075" heatid="4908" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4286" nation="GER" region="02" clubid="3328" name="SC DELPHIN Ingolstadt">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Rafaela" gender="F" lastname="Averbeck" nation="GER" license="295302" athleteid="3332">
              <RESULTS>
                <RESULT eventid="1059" points="513" swimtime="00:01:03.59" resultid="3333" heatid="4665" lane="2" entrytime="00:01:03.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="564" swimtime="00:04:43.74" resultid="3334" heatid="4762" lane="4" entrytime="00:04:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="100" swimtime="00:01:07.71" />
                    <SPLIT distance="150" swimtime="00:01:44.17" />
                    <SPLIT distance="200" swimtime="00:02:20.46" />
                    <SPLIT distance="250" swimtime="00:02:56.91" />
                    <SPLIT distance="300" swimtime="00:03:33.13" />
                    <SPLIT distance="350" swimtime="00:04:09.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:14.00" eventid="1978" heatid="4834" lane="3" />
                <ENTRY entrytime="00:09:56.68" eventid="2020" heatid="4875" lane="1">
                  <MEETINFO qualificationtime="00:09:56.68" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Daniel" gender="M" lastname="Chen" nation="GER" license="280055" athleteid="3338">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.60" eventid="1971" heatid="4817" lane="5" />
                <ENTRY entrytime="00:01:06.40" eventid="2013" heatid="4869" lane="1" />
                <ENTRY entrytime="00:00:28.40" eventid="2103" heatid="4941" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Jonas" gender="M" lastname="Drieling" nation="GER" license="280053" athleteid="3345">
              <RESULTS>
                <RESULT eventid="1778" points="518" swimtime="00:01:00.29" resultid="3346" heatid="4713" lane="2" entrytime="00:01:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="522" swimtime="00:00:27.59" resultid="3347" heatid="4742" lane="5" entrytime="00:00:28.40" />
                <RESULT eventid="1834" points="542" swimtime="00:00:24.84" resultid="3348" heatid="4771" lane="2" entrytime="00:00:25.60" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.40" eventid="1971" heatid="4822" lane="1" />
                <ENTRY entrytime="00:01:03.40" eventid="2027" heatid="4880" lane="6" />
                <ENTRY entrytime="00:00:26.90" eventid="2103" heatid="4945" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Olivia" gender="F" lastname="Gerrard" nation="GER" license="266868" athleteid="3352">
              <RESULTS>
                <RESULT eventid="1059" points="555" swimtime="00:01:01.93" resultid="3353" heatid="4669" lane="2" entrytime="00:01:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="531" swimtime="00:01:07.93" resultid="3354" heatid="4722" lane="1" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="547" swimtime="00:00:29.80" resultid="3355" heatid="4800" lane="1" entrytime="00:00:29.80" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:08.80" eventid="2006" heatid="4864" lane="4" />
                <ENTRY entrytime="00:02:31.20" eventid="2055" heatid="4904" lane="6" />
                <ENTRY entrytime="00:02:26.80" eventid="2096" heatid="4937" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Simon" gender="M" lastname="Göpffarth" nation="GER" license="316788" athleteid="3359">
              <RESULTS>
                <RESULT eventid="1749" points="455" swimtime="00:02:09.18" resultid="3360" heatid="4677" lane="5" entrytime="00:02:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                    <SPLIT distance="100" swimtime="00:01:02.55" />
                    <SPLIT distance="150" swimtime="00:01:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="440" swimtime="00:00:26.63" resultid="3361" heatid="4767" lane="5" entrytime="00:00:26.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Fabian" gender="M" lastname="Heinemann" nation="GER" license="313851" athleteid="3362">
              <RESULTS>
                <RESULT eventid="1778" points="444" swimtime="00:01:03.45" resultid="3363" heatid="4710" lane="6" entrytime="00:01:03.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="436" swimtime="00:00:29.30" resultid="3364" heatid="4740" lane="6" entrytime="00:00:30.00" />
                <RESULT eventid="1834" points="518" swimtime="00:00:25.22" resultid="3365" heatid="4770" lane="6" entrytime="00:00:26.00" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.40" eventid="1971" heatid="4820" lane="2" />
                <ENTRY entrytime="00:01:04.20" eventid="2027" heatid="4878" lane="2" />
                <ENTRY entrytime="00:00:28.00" eventid="2103" heatid="4942" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Larissa" gender="F" lastname="Heinemann" nation="GER" license="313844" athleteid="3369">
              <RESULTS>
                <RESULT eventid="1059" points="540" swimtime="00:01:02.48" resultid="3370" heatid="4667" lane="1" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="487" swimtime="00:01:12.02" resultid="3371" heatid="4733" lane="3" entrytime="00:01:11.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="483" swimtime="00:00:31.06" resultid="3372" heatid="4795" lane="3" entrytime="00:00:31.60" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:19.90" eventid="1992" heatid="4852" lane="1" />
                <ENTRY entrytime="00:00:28.40" eventid="2082" heatid="4920" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Joshua" gender="M" lastname="Hollweck" nation="GER" license="313850" athleteid="3375">
              <RESULTS>
                <RESULT eventid="1778" points="506" swimtime="00:01:00.76" resultid="3376" heatid="4712" lane="3" entrytime="00:01:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="521" swimtime="00:02:16.24" resultid="3377" heatid="4753" lane="1" entrytime="00:02:15.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:04.45" />
                    <SPLIT distance="150" swimtime="00:01:46.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.20" eventid="1971" heatid="4822" lane="2" />
                <ENTRY entrytime="00:02:16.40" eventid="2041" heatid="4893" lane="1" />
                <ENTRY entrytime="00:00:28.10" eventid="2103" heatid="4942" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Iberle" nation="GER" license="313842" athleteid="3381">
              <RESULTS>
                <RESULT eventid="1059" points="482" swimtime="00:01:04.89" resultid="3382" heatid="4664" lane="6" entrytime="00:01:04.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="535" swimtime="00:04:48.71" resultid="3383" heatid="4759" lane="3" entrytime="00:04:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:46.30" />
                    <SPLIT distance="200" swimtime="00:02:23.26" />
                    <SPLIT distance="250" swimtime="00:02:59.97" />
                    <SPLIT distance="300" swimtime="00:03:36.96" />
                    <SPLIT distance="350" swimtime="00:04:13.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:20.80" eventid="1978" heatid="4829" lane="4" />
                <ENTRY entrytime="00:02:38.20" eventid="2055" heatid="4898" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lina" gender="F" lastname="Kapfer" nation="GER" license="322567" athleteid="3386">
              <RESULTS>
                <RESULT eventid="1799" points="460" swimtime="00:01:13.39" resultid="3387" heatid="4729" lane="1" entrytime="00:01:14.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="458" swimtime="00:02:54.52" resultid="3388" heatid="4780" lane="1" entrytime="00:02:54.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:08.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Maria" gender="F" lastname="Kapfer" nation="GER" license="322566" athleteid="3389">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.90" eventid="2034" heatid="4884" lane="4" />
                <ENTRY entrytime="00:02:36.40" eventid="2096" heatid="4932" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sara Maria" gender="F" lastname="Krönert" nation="GER" license="339853" athleteid="3392">
              <ENTRIES>
                <ENTRY entrytime="00:02:33.80" eventid="2096" heatid="4933" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Kuhls" nation="GER" license="265730" athleteid="3394">
              <RESULTS>
                <RESULT eventid="1059" points="540" swimtime="00:01:02.49" resultid="3395" heatid="4668" lane="3" entrytime="00:01:02.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="519" swimtime="00:04:51.65" resultid="3396" heatid="4760" lane="5" entrytime="00:04:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.65" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:46.16" />
                    <SPLIT distance="200" swimtime="00:02:23.54" />
                    <SPLIT distance="250" swimtime="00:03:01.38" />
                    <SPLIT distance="300" swimtime="00:03:38.73" />
                    <SPLIT distance="350" swimtime="00:04:16.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:17.60" eventid="1978" heatid="4832" lane="5" />
                <ENTRY entrytime="00:00:33.40" eventid="2034" heatid="4885" lane="4" />
                <ENTRY entrytime="00:00:28.60" eventid="2082" heatid="4918" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lukas" gender="M" lastname="Meilinger" nation="GER" license="246338" athleteid="3400">
              <RESULTS>
                <RESULT eventid="1834" points="490" swimtime="00:00:25.69" resultid="3401" heatid="4771" lane="4" entrytime="00:00:25.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Raphael" gender="M" lastname="Mooser" nation="GER" license="280056" athleteid="3402">
              <RESULTS>
                <RESULT eventid="1763" points="450" swimtime="00:01:12.52" resultid="3403" heatid="4699" lane="1" entrytime="00:01:10.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="436" swimtime="00:02:24.53" resultid="3404" heatid="4750" lane="4" entrytime="00:02:23.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:09.64" />
                    <SPLIT distance="150" swimtime="00:01:50.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.80" eventid="1985" heatid="4842" lane="4" />
                <ENTRY entrytime="00:02:31.20" eventid="2089" heatid="4928" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Sascha" gender="M" lastname="Santa" nation="GER" license="279042" athleteid="3407">
              <RESULTS>
                <RESULT eventid="1749" points="573" swimtime="00:01:59.60" resultid="3408" heatid="4682" lane="5" entrytime="00:02:00.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                    <SPLIT distance="100" swimtime="00:00:58.52" />
                    <SPLIT distance="150" swimtime="00:01:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="486" swimtime="00:02:19.36" resultid="3409" heatid="4751" lane="3" entrytime="00:02:21.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="100" swimtime="00:01:06.83" />
                    <SPLIT distance="150" swimtime="00:01:47.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.60" eventid="1971" heatid="4821" lane="2" />
                <ENTRY entrytime="00:04:13.80" eventid="2075" heatid="4910" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Johanna" gender="F" lastname="Schmid" nation="GER" license="266871" athleteid="3412">
              <RESULTS>
                <RESULT eventid="1756" points="547" swimtime="00:00:35.20" resultid="3413" heatid="4691" lane="5" entrytime="00:00:35.60" />
                <RESULT eventid="1799" points="506" swimtime="00:01:11.10" resultid="3414" heatid="4735" lane="6" entrytime="00:01:11.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="478" swimtime="00:02:52.00" resultid="3415" heatid="4781" lane="5" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:07.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:18.90" eventid="1992" heatid="4853" lane="6" />
                <ENTRY entrytime="00:02:35.40" eventid="2055" heatid="4900" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Vanessa" gender="F" lastname="Waal" nation="GER" license="301334" athleteid="3418">
              <RESULTS>
                <RESULT eventid="1059" points="503" swimtime="00:01:04.00" resultid="3419" heatid="4666" lane="1" entrytime="00:01:03.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="480" swimtime="00:01:12.35" resultid="3420" heatid="4731" lane="5" entrytime="00:01:12.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:20.50" eventid="1978" heatid="4830" lane="5" />
                <ENTRY entrytime="00:00:29.40" eventid="2082" heatid="4915" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4292" nation="GER" region="02" clubid="4087" name="SC Prinz Eugen München">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Alexander Philip" gender="M" lastname="Adami" nation="GER" license="297199" swrid="4829107" athleteid="4103">
              <RESULTS>
                <RESULT eventid="1778" points="441" swimtime="00:01:03.60" resultid="4104" heatid="4710" lane="2" entrytime="00:01:03.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.07" eventid="1971" heatid="4816" lane="6" />
                <ENTRY entrytime="00:00:28.11" eventid="2103" heatid="4941" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Juliana Andrea" gender="F" lastname="Adami" nation="GER" license="297636" swrid="4829108" athleteid="4107">
              <RESULTS>
                <RESULT eventid="1059" points="522" swimtime="00:01:03.22" resultid="4108" heatid="4666" lane="4" entrytime="00:01:03.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="509" swimtime="00:01:10.94" resultid="4109" heatid="4730" lane="2" entrytime="00:01:13.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="485" swimtime="00:00:31.02" resultid="4110" heatid="4798" lane="3" entrytime="00:00:30.72" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:19.76" eventid="1978" heatid="4831" lane="6" />
                <ENTRY entrytime="00:01:09.83" eventid="2006" heatid="4864" lane="2" />
                <ENTRY entrytime="00:02:36.27" eventid="2055" heatid="4899" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Lyubomir" gender="M" lastname="Agov" nation="GER" license="372659" athleteid="4114">
              <RESULTS>
                <RESULT eventid="1763" points="693" swimtime="00:01:02.84" resultid="4115" heatid="4701" lane="3" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1884" points="702" swimtime="00:01:02.55" resultid="5357" heatid="4704" lane="4" entrytime="00:01:02.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:26.95" eventid="1985" heatid="4848" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Markus" gender="M" lastname="Fischer" nation="GER" license="297634" athleteid="4117">
              <RESULTS>
                <RESULT eventid="1749" points="520" swimtime="00:02:03.55" resultid="4118" heatid="4681" lane="1" entrytime="00:02:02.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                    <SPLIT distance="100" swimtime="00:00:59.44" />
                    <SPLIT distance="150" swimtime="00:01:31.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="468" swimtime="00:02:16.01" resultid="4119" heatid="4790" lane="5" entrytime="00:02:13.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="150" swimtime="00:01:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="479" swimtime="00:02:14.99" resultid="5500" heatid="5504" lane="2" entrytime="00:02:16.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                    <SPLIT distance="150" swimtime="00:01:40.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.86" eventid="1971" heatid="4819" lane="1" />
                <ENTRY entrytime="00:01:02.22" eventid="2013" heatid="4871" lane="1" />
                <ENTRY entrytime="00:04:22.05" eventid="2075" heatid="4909" lane="2" />
                <ENTRY entrytime="00:09:07.54" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:07.54" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Jasper" gender="M" lastname="Glindemann" nation="GER" license="309671" athleteid="4124">
              <RESULTS>
                <RESULT eventid="1763" points="510" swimtime="00:01:09.57" resultid="4125" heatid="4698" lane="5" entrytime="00:01:10.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="446" swimtime="00:02:23.40" resultid="4126" heatid="4749" lane="4" entrytime="00:02:27.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                    <SPLIT distance="100" swimtime="00:01:09.47" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.10" eventid="1985" heatid="4845" lane="5" />
                <ENTRY entrytime="00:01:08.56" eventid="2027" heatid="4877" lane="2" />
                <ENTRY entrytime="00:02:36.40" eventid="2089" heatid="4927" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Kevin" gender="M" lastname="Hültner" nation="GER" license="250305" athleteid="4130">
              <RESULTS>
                <RESULT eventid="1763" points="544" swimtime="00:01:08.11" resultid="4131" heatid="4701" lane="6" entrytime="00:01:06.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.56" eventid="1985" heatid="4847" lane="6" />
                <ENTRY entrytime="00:02:31.29" eventid="2089" heatid="4927" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Laura" gender="F" lastname="Jaeschke" nation="GER" license="326712" athleteid="4134">
              <RESULTS>
                <RESULT eventid="1059" points="447" swimtime="00:01:06.55" resultid="4135" heatid="4663" lane="6" entrytime="00:01:04.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="537" swimtime="00:04:48.37" resultid="4136" heatid="4759" lane="5" entrytime="00:04:54.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:01:45.87" />
                    <SPLIT distance="200" swimtime="00:02:22.36" />
                    <SPLIT distance="250" swimtime="00:02:59.13" />
                    <SPLIT distance="300" swimtime="00:03:36.30" />
                    <SPLIT distance="350" swimtime="00:04:13.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Patryk" gender="M" lastname="Laszyca" nation="GER" license="290977" athleteid="4137">
              <RESULTS>
                <RESULT eventid="1778" points="522" swimtime="00:01:00.13" resultid="4138" heatid="4716" lane="1" entrytime="00:00:59.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="547" swimtime="00:00:24.76" resultid="4139" heatid="4774" lane="1" entrytime="00:00:24.93" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.86" eventid="1971" heatid="4824" lane="4" />
                <ENTRY entrytime="00:01:03.35" eventid="2027" heatid="4881" lane="6" />
                <ENTRY entrytime="00:00:27.31" eventid="2103" heatid="4944" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Hanna" gender="F" lastname="Pfannes" nation="GER" license="301469" athleteid="4143">
              <RESULTS>
                <RESULT eventid="1756" points="495" swimtime="00:00:36.40" resultid="4144" heatid="4689" lane="6" entrytime="00:00:37.09" />
                <RESULT eventid="1841" points="525" swimtime="00:02:46.80" resultid="4145" heatid="4783" lane="5" entrytime="00:02:45.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:18.36" />
                    <SPLIT distance="150" swimtime="00:02:01.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:16.20" eventid="1992" heatid="4857" lane="1" />
                <ENTRY entrytime="00:00:33.82" eventid="2034" heatid="4884" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Amelie" gender="F" lastname="Zachenhuber" nation="GER" license="304970" athleteid="4148">
              <RESULTS>
                <RESULT eventid="1059" points="593" swimtime="00:01:00.57" resultid="4149" heatid="4671" lane="2" entrytime="00:01:01.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="554" swimtime="00:00:35.05" resultid="4150" heatid="4692" lane="5" entrytime="00:00:34.57" />
                <RESULT eventid="1785" points="503" swimtime="00:01:09.18" resultid="4151" heatid="4722" lane="6" entrytime="00:01:08.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="508" swimtime="00:01:11.02" resultid="4152" heatid="4734" lane="5" entrytime="00:01:10.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="548" swimtime="00:00:29.79" resultid="4153" heatid="4961" lane="2" entrytime="00:00:29.32" />
                <RESULT eventid="1940" points="600" swimtime="00:00:28.89" resultid="5513" heatid="5517" lane="2" entrytime="00:00:29.79" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:16.36" eventid="1992" heatid="4857" lane="6" />
                <ENTRY entrytime="00:01:07.60" eventid="2006" heatid="4865" lane="1" />
                <ENTRY entrytime="00:00:31.85" eventid="2034" heatid="4889" lane="6" />
                <ENTRY entrytime="00:00:27.53" eventid="2082" heatid="4922" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="570" swimtime="00:01:49.11" resultid="4158" heatid="4805" lane="3" entrytime="00:01:53.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="100" swimtime="00:00:56.68" />
                    <SPLIT distance="150" swimtime="00:01:24.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4117" number="1" />
                    <RELAYPOSITION athleteid="4114" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4103" number="3" reactiontime="+47" />
                    <RELAYPOSITION athleteid="4137" number="4" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6524" nation="GER" region="02" clubid="2699" name="SC Regensburg">
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Julia Maria" gender="F" lastname="Grasser" nation="GER" license="179987" athleteid="2700">
              <RESULTS>
                <RESULT eventid="1813" points="495" swimtime="00:02:31.17" resultid="2701" heatid="4746" lane="5" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:11.04" />
                    <SPLIT distance="150" swimtime="00:01:51.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:14.15" eventid="1978" heatid="4834" lane="4" />
                <ENTRY entrytime="00:01:07.16" eventid="2006" heatid="4867" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Maximilian" gender="M" lastname="Peter" nation="GER" license="228199" athleteid="2704">
              <RESULTS>
                <RESULT eventid="1806" points="414" swimtime="00:00:29.81" resultid="2705" heatid="4740" lane="4" entrytime="00:00:29.30" />
                <RESULT eventid="1848" points="454" swimtime="00:02:17.40" resultid="2706" heatid="4791" lane="5" entrytime="00:02:13.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:42.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:02.14" eventid="2013" heatid="4872" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4296" nation="GER" region="02" clubid="3640" name="SC Wfr. München">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Marvin" gender="M" lastname="Christmann" nation="GER" license="248439" athleteid="3656">
              <RESULTS>
                <RESULT eventid="1763" points="464" swimtime="00:01:11.82" resultid="3657" heatid="4699" lane="5" entrytime="00:01:10.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="498" swimtime="00:00:25.56" resultid="3658" heatid="4773" lane="6" entrytime="00:00:25.13" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.36" eventid="1985" heatid="4844" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Dominic" gender="M" lastname="Ehinlanwo" nation="GER" license="302032" athleteid="3660">
              <RESULTS>
                <RESULT eventid="1749" points="583" swimtime="00:01:58.92" resultid="3661" heatid="4684" lane="6" entrytime="00:01:57.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                    <SPLIT distance="100" swimtime="00:00:56.89" />
                    <SPLIT distance="150" swimtime="00:01:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="549" swimtime="00:00:24.73" resultid="3662" heatid="4773" lane="2" entrytime="00:00:25.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Bruno" gender="M" lastname="Hediger" nation="GER" license="387694" athleteid="3663">
              <RESULTS>
                <RESULT eventid="1778" points="579" swimtime="00:00:58.10" resultid="3664" heatid="4714" lane="5" entrytime="00:00:59.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="601" swimtime="00:02:09.84" resultid="3665" heatid="4754" lane="1" entrytime="00:02:11.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                    <SPLIT distance="150" swimtime="00:01:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1898" points="585" swimtime="00:00:57.90" resultid="5458" heatid="4717" lane="6" entrytime="00:00:58.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julius" gender="M" lastname="Hirschberg" nation="GER" license="333024" athleteid="3666">
              <RESULTS>
                <RESULT eventid="1778" points="467" swimtime="00:01:02.41" resultid="3667" heatid="4711" lane="3" entrytime="00:01:02.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="514" swimtime="00:00:25.28" resultid="3668" heatid="4771" lane="6" entrytime="00:00:25.73" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:27.26" eventid="2103" heatid="4944" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Matthias" gender="M" lastname="Killiches" nation="GER" license="73649" athleteid="3670">
              <RESULTS>
                <RESULT eventid="1763" points="535" swimtime="00:01:08.50" resultid="3671" heatid="4700" lane="3" entrytime="00:01:07.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.09" eventid="1985" heatid="4845" lane="2" />
                <ENTRY entrytime="00:02:28.00" eventid="2089" heatid="4930" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Jörg" gender="M" lastname="Lukashov" nation="GER" license="252298" athleteid="3674">
              <RESULTS>
                <RESULT eventid="1763" points="593" swimtime="00:01:06.19" resultid="3675" heatid="4702" lane="1" entrytime="00:01:05.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="605" swimtime="00:00:23.95" resultid="3676" heatid="4777" lane="1" entrytime="00:00:24.05" />
                <RESULT eventid="1947" points="599" swimtime="00:00:24.03" resultid="5471" heatid="4778" lane="6" entrytime="00:00:23.95" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.22" eventid="1971" heatid="4825" lane="5" />
                <ENTRY entrytime="00:00:59.00" eventid="2027" heatid="4879" lane="4" />
                <ENTRY entrytime="00:00:25.82" eventid="2103" heatid="4946" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Frida" gender="F" lastname="Mayr" nation="GER" license="356519" athleteid="3680">
              <RESULTS>
                <RESULT eventid="1059" points="476" swimtime="00:01:05.16" resultid="3681" heatid="4668" lane="1" entrytime="00:01:02.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="452" swimtime="00:00:31.76" resultid="3682" heatid="4795" lane="4" entrytime="00:00:31.62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Viola Jasmine" gender="F" lastname="Provost" nation="GER" license="329228" athleteid="3683">
              <RESULTS>
                <RESULT eventid="1059" points="545" swimtime="00:01:02.32" resultid="3684" heatid="4669" lane="1" entrytime="00:01:02.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:28.24" eventid="2082" heatid="4921" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Roman" gender="M" lastname="Roelen" nation="GER" license="283816" athleteid="3686">
              <RESULTS>
                <RESULT eventid="1749" points="443" swimtime="00:02:10.28" resultid="3687" heatid="4676" lane="4" entrytime="00:02:11.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:03.31" />
                    <SPLIT distance="150" swimtime="00:01:37.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1971" heatid="4813" lane="4" />
                <ENTRY entrytime="00:04:38.00" eventid="2075" heatid="4907" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Alexander" gender="M" lastname="Roschlaub" nation="GER" license="140735" athleteid="3690">
              <RESULTS>
                <RESULT eventid="1749" points="598" swimtime="00:01:57.91" resultid="3691" heatid="4682" lane="4" entrytime="00:02:00.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="100" swimtime="00:00:57.55" />
                    <SPLIT distance="150" swimtime="00:01:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="585" swimtime="00:00:24.22" resultid="3692" heatid="4775" lane="1" entrytime="00:00:24.50" />
                <RESULT eventid="1947" points="607" swimtime="00:00:23.92" resultid="5475" heatid="5478" lane="5" entrytime="00:00:24.22" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.31" eventid="1971" heatid="4827" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Alexandra" gender="F" lastname="Schäffler" nation="GER" license="231075" athleteid="3694">
              <RESULTS>
                <RESULT eventid="1756" points="484" swimtime="00:00:36.68" resultid="3695" heatid="4691" lane="6" entrytime="00:00:35.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Manuel" gender="M" lastname="Straßl" nation="GER" license="132560" athleteid="3696">
              <RESULTS>
                <RESULT eventid="1806" points="479" swimtime="00:00:28.38" resultid="3697" heatid="4743" lane="5" entrytime="00:00:28.23" />
                <RESULT eventid="1834" points="595" swimtime="00:00:24.08" resultid="3698" heatid="4774" lane="4" entrytime="00:00:24.70" />
                <RESULT eventid="1947" points="585" swimtime="00:00:24.22" resultid="5473" heatid="5478" lane="4" entrytime="00:00:24.08" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.67" eventid="1971" heatid="4823" lane="1" />
                <ENTRY entrytime="00:01:03.02" eventid="2027" heatid="4880" lane="1" />
                <ENTRY entrytime="00:00:27.00" eventid="2103" heatid="4946" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="570" swimtime="00:01:49.13" resultid="3702" heatid="4805" lane="5" entrytime="00:02:00.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:00:59.36" />
                    <SPLIT distance="150" swimtime="00:01:25.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3696" number="1" />
                    <RELAYPOSITION athleteid="3670" number="2" reactiontime="+19" />
                    <RELAYPOSITION athleteid="3663" number="3" reactiontime="+18" />
                    <RELAYPOSITION athleteid="3674" number="4" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="(Zeit: 19:29), Der 3. Schwimmer verließ den Startblock bevor der 2. Schwimmer angeschlagen hat." eventid="2048" status="DSQ" swimtime="00:01:51.46" resultid="3704" heatid="4805" lane="1" entrytime="00:02:02.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                    <SPLIT distance="100" swimtime="00:01:00.81" />
                    <SPLIT distance="150" swimtime="00:01:27.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3690" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3656" number="2" reactiontime="+39" status="DSQ" />
                    <RELAYPOSITION athleteid="3666" number="3" reactiontime="+33" status="DSQ" />
                    <RELAYPOSITION athleteid="3660" number="4" reactiontime="+43" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:42.63" eventid="2232" heatid="4811" lane="4" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4344" nation="GER" region="02" clubid="3263" name="SCHWIMMVEREIN AUGSBURG 1911 e.V." shortname="SCHWIMMVEREIN AUGSBURG 1911 e.">
          <ATHLETES>
            <ATHLETE birthdate="1989-01-01" firstname="Nadine" gender="F" lastname="Bender" nation="GER" license="197915" athleteid="3264">
              <RESULTS>
                <RESULT eventid="1059" points="619" swimtime="00:00:59.71" resultid="3265" heatid="4673" lane="4" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="543" swimtime="00:01:07.45" resultid="3266" heatid="4723" lane="2" entrytime="00:01:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="630" swimtime="00:00:59.36" resultid="5325" heatid="5317" lane="4" entrytime="00:00:59.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1891" points="563" swimtime="00:01:06.64" resultid="5390" heatid="5391" lane="6" entrytime="00:01:07.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:08.50" eventid="1978" heatid="4837" lane="2" />
                <ENTRY entrytime="00:00:30.60" eventid="2034" heatid="4888" lane="4" />
                <ENTRY entrytime="00:00:27.30" eventid="2082" heatid="4922" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Cara" gender="F" lastname="Gallina" nation="GER" license="299199" athleteid="3270">
              <RESULTS>
                <RESULT eventid="1059" points="556" swimtime="00:01:01.90" resultid="3271" heatid="4664" lane="3" entrytime="00:01:03.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="522" swimtime="00:00:30.26" resultid="3272" heatid="4796" lane="1" entrytime="00:00:31.50" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:16.00" eventid="1978" heatid="4833" lane="6" />
                <ENTRY entrytime="00:00:28.51" eventid="2082" heatid="4919" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Matthias" gender="M" lastname="Kopfmüller" nation="GER" license="137031" athleteid="3275">
              <RESULTS>
                <RESULT eventid="1778" points="545" swimtime="00:00:59.28" resultid="3276" heatid="4715" lane="2" entrytime="00:00:58.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="582" swimtime="00:00:24.26" resultid="3277" heatid="4775" lane="4" entrytime="00:00:23.40" />
                <RESULT eventid="5443" points="573" swimtime="00:00:24.39" resultid="5450" heatid="5452" lane="3" entrytime="00:00:24.26" />
                <RESULT eventid="1947" points="601" swimtime="00:00:24.00" resultid="5477" heatid="5478" lane="6" entrytime="00:00:24.26" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:51.90" eventid="1971" heatid="4827" lane="2" />
                <ENTRY entrytime="00:00:25.90" eventid="2103" heatid="4945" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Andreas" gender="M" lastname="Kornes" nation="GER" license="075398" athleteid="3280">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.40" eventid="1985" heatid="4846" lane="4" />
                <ENTRY entrytime="00:02:23.50" eventid="2089" heatid="4928" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Michelle" gender="F" lastname="Lienhart" nation="GER" license="203026" athleteid="3283">
              <RESULTS>
                <RESULT eventid="1059" points="626" swimtime="00:00:59.49" resultid="3284" heatid="4672" lane="4" entrytime="00:00:58.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="553" swimtime="00:01:09.01" resultid="3285" heatid="4734" lane="3" entrytime="00:01:06.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="573" swimtime="00:00:29.35" resultid="3286" heatid="4800" lane="2" entrytime="00:00:29.44" />
                <RESULT eventid="1863" points="625" swimtime="00:00:59.52" resultid="5322" heatid="4675" lane="1" entrytime="00:00:59.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="569" swimtime="00:00:29.41" resultid="5510" heatid="4802" lane="6" entrytime="00:00:29.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Oliver" gender="M" lastname="Lienhart" nation="GER" license="248518" athleteid="3287">
              <RESULTS>
                <RESULT eventid="1763" points="480" swimtime="00:01:10.98" resultid="3288" heatid="4699" lane="6" entrytime="00:01:10.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="427" swimtime="00:02:20.25" resultid="3289" heatid="4788" lane="6" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:08.15" />
                    <SPLIT distance="150" swimtime="00:01:44.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.74" eventid="1971" heatid="4817" lane="6" />
                <ENTRY entrytime="00:01:03.68" eventid="2027" heatid="4878" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Leonie" gender="F" lastname="Mathe" nation="GER" license="215384" athleteid="3292">
              <RESULTS>
                <RESULT eventid="1059" points="624" swimtime="00:00:59.56" resultid="3293" heatid="4674" lane="5" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="609" swimtime="00:00:33.96" resultid="3294" heatid="4692" lane="2" entrytime="00:00:34.00" />
                <RESULT eventid="1841" points="551" swimtime="00:02:44.09" resultid="3295" heatid="4784" lane="6" entrytime="00:02:47.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:19.46" />
                    <SPLIT distance="150" swimtime="00:02:02.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1877" points="649" swimtime="00:00:33.26" resultid="5348" heatid="4695" lane="6" entrytime="00:00:33.96" />
                <RESULT eventid="1954" points="586" swimtime="00:02:40.74" resultid="5487" heatid="5491" lane="2" entrytime="00:02:44.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:02:00.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:15.50" eventid="1992" heatid="4855" lane="2" />
                <ENTRY entrytime="00:00:27.50" eventid="2082" heatid="4923" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Laura" gender="F" lastname="Popp" nation="GER" license="178550" athleteid="3298">
              <RESULTS>
                <RESULT eventid="1756" points="588" swimtime="00:00:34.36" resultid="3299" heatid="4694" lane="2" entrytime="00:00:33.60" />
                <RESULT eventid="1799" points="532" swimtime="00:01:09.92" resultid="3300" heatid="4735" lane="2" entrytime="00:01:07.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="588" swimtime="00:02:40.61" resultid="3301" heatid="4782" lane="3" entrytime="00:02:38.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:17.35" />
                    <SPLIT distance="150" swimtime="00:01:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1877" points="609" swimtime="00:00:33.97" resultid="5352" heatid="5355" lane="5" entrytime="00:00:34.36" />
                <RESULT eventid="1919" points="537" swimtime="00:01:09.69" resultid="5398" heatid="5404" lane="3" entrytime="00:01:09.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1954" points="589" swimtime="00:02:40.46" resultid="5484" heatid="4785" lane="6" entrytime="00:02:40.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="100" swimtime="00:01:17.14" />
                    <SPLIT distance="150" swimtime="00:01:58.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:12.90" eventid="1992" heatid="4857" lane="4" />
                <ENTRY entrytime="00:02:27.30" eventid="2055" heatid="4902" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Lea" gender="F" lastname="Preußner" nation="GER" license="282176" athleteid="3304">
              <RESULTS>
                <RESULT eventid="1771" points="456" swimtime="00:05:36.85" resultid="3305" heatid="4707" lane="2" entrytime="00:05:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                    <SPLIT distance="100" swimtime="00:01:15.06" />
                    <SPLIT distance="150" swimtime="00:01:57.70" />
                    <SPLIT distance="200" swimtime="00:02:39.90" />
                    <SPLIT distance="250" swimtime="00:03:28.09" />
                    <SPLIT distance="300" swimtime="00:04:19.03" />
                    <SPLIT distance="350" swimtime="00:04:58.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="426" swimtime="00:01:15.31" resultid="3306" heatid="4731" lane="2" entrytime="00:01:12.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Paul" gender="M" lastname="Pucknus" nation="GER" license="264470" athleteid="3307">
              <RESULTS>
                <RESULT eventid="1778" points="486" swimtime="00:01:01.58" resultid="3308" heatid="4711" lane="2" entrytime="00:01:02.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="406" swimtime="00:02:22.55" resultid="3309" heatid="4787" lane="6" entrytime="00:02:22.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:46.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.65" eventid="1971" heatid="4815" lane="1" />
                <ENTRY entrytime="00:02:17.06" eventid="2041" heatid="4894" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Matthias" gender="M" lastname="Schwab" nation="GER" license="132395" athleteid="3312">
              <RESULTS>
                <RESULT eventid="1778" points="551" swimtime="00:00:59.07" resultid="3313" heatid="4715" lane="1" entrytime="00:00:59.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1898" points="555" swimtime="00:00:58.94" resultid="5463" heatid="5465" lane="1" entrytime="00:00:59.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.20" eventid="1985" heatid="4847" lane="1" />
                <ENTRY entrytime="00:00:25.50" eventid="2103" heatid="4947" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Denis" gender="M" lastname="Sczesny" nation="GER" license="350186" athleteid="3316">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.67" eventid="1985" heatid="4841" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Oliver" gender="M" lastname="Sczesny" nation="GER" license="330650" athleteid="3318">
              <RESULTS>
                <RESULT eventid="1763" points="646" swimtime="00:01:04.32" resultid="3319" heatid="4702" lane="5" entrytime="00:01:04.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1884" points="660" swimtime="00:01:03.87" resultid="5363" heatid="5368" lane="4" entrytime="00:01:04.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.26" eventid="1985" heatid="4846" lane="1" />
                <ENTRY entrytime="00:02:23.53" eventid="2089" heatid="4930" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Mark" gender="M" lastname="Toprak" nation="GER" license="346434" athleteid="3322">
              <RESULTS>
                <RESULT eventid="1749" points="526" swimtime="00:02:03.09" resultid="3323" heatid="4680" lane="5" entrytime="00:02:03.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="100" swimtime="00:00:59.92" />
                    <SPLIT distance="150" swimtime="00:01:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="425" swimtime="00:01:04.38" resultid="3324" heatid="4710" lane="4" entrytime="00:01:02.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.57" eventid="1971" heatid="4820" lane="1" />
                <ENTRY entrytime="00:02:34.84" eventid="2089" heatid="4927" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="2062" points="596" swimtime="00:02:03.58" resultid="3327" heatid="4807" lane="5" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:36.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3264" number="1" />
                    <RELAYPOSITION athleteid="3298" number="2" />
                    <RELAYPOSITION athleteid="3283" number="3" />
                    <RELAYPOSITION athleteid="3292" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6399" nation="GER" region="02" clubid="3208" name="SG - Elsenfeld/Kleinwallstadt">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Stefanie" gender="F" lastname="Göller" nation="GER" license="245438" athleteid="3217">
              <RESULTS>
                <RESULT eventid="1059" points="570" swimtime="00:01:01.39" resultid="3218" heatid="4668" lane="6" entrytime="00:01:02.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="461" swimtime="00:01:11.21" resultid="3219" heatid="4720" lane="6" entrytime="00:01:11.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="478" swimtime="00:01:12.45" resultid="3220" heatid="4731" lane="3" entrytime="00:01:12.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="474" swimtime="00:00:31.25" resultid="3221" heatid="4796" lane="5" entrytime="00:00:31.42" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:33.48" eventid="2034" heatid="4885" lane="5" />
                <ENTRY entrytime="00:00:28.76" eventid="2082" heatid="4918" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Noelle" gender="F" lastname="Ronalter" nation="GER" license="288664" athleteid="3224">
              <RESULTS>
                <RESULT eventid="1059" points="484" swimtime="00:01:04.80" resultid="3225" heatid="4662" lane="2" entrytime="00:01:05.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="391" swimtime="00:01:15.23" resultid="3226" heatid="4718" lane="3" entrytime="00:01:13.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="400" swimtime="00:01:16.87" resultid="3227" heatid="4728" lane="2" entrytime="00:01:15.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:34.21" eventid="2034" heatid="4883" lane="3" />
                <ENTRY entrytime="00:00:29.91" eventid="2082" heatid="4914" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5085" nation="GER" region="02" clubid="4172" name="SG Bamberg">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Benedikt" gender="M" lastname="Dörfler" nation="GER" license="169778" athleteid="4173">
              <RESULTS>
                <RESULT eventid="1749" points="487" swimtime="00:02:06.25" resultid="4174" heatid="4680" lane="1" entrytime="00:02:03.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:01:00.07" />
                    <SPLIT distance="150" swimtime="00:01:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="420" swimtime="00:00:29.67" resultid="4175" heatid="4740" lane="3" entrytime="00:00:29.26" />
                <RESULT eventid="1848" points="466" swimtime="00:02:16.16" resultid="4176" heatid="4788" lane="4" entrytime="00:02:18.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:06.38" />
                    <SPLIT distance="150" swimtime="00:01:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="459" swimtime="00:02:16.91" resultid="5502" heatid="5504" lane="1" entrytime="00:02:16.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:41.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.76" eventid="1971" heatid="4819" lane="5" />
                <ENTRY entrytime="00:01:01.77" eventid="2013" heatid="4871" lane="5" />
                <ENTRY entrytime="00:04:23.39" eventid="2075" heatid="4909" lane="1" />
                <ENTRY entrytime="00:00:28.86" eventid="2103" heatid="4940" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Nikolas" gender="M" lastname="Häfner" nation="GER" license="196438" athleteid="4181">
              <RESULTS>
                <RESULT eventid="1806" points="536" swimtime="00:00:27.35" resultid="4182" heatid="4741" lane="3" entrytime="00:00:26.55" />
                <RESULT eventid="1834" points="529" swimtime="00:00:25.05" resultid="4183" heatid="4773" lane="1" entrytime="00:00:25.03" />
                <RESULT eventid="1848" points="514" swimtime="00:02:11.82" resultid="4184" heatid="4791" lane="3" entrytime="00:02:05.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:02.80" />
                    <SPLIT distance="150" swimtime="00:01:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1912" points="553" swimtime="00:00:27.06" resultid="5408" heatid="4744" lane="5" entrytime="00:00:27.35" />
                <RESULT eventid="1961" points="522" swimtime="00:02:11.18" resultid="5495" heatid="4792" lane="5" entrytime="00:02:11.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:03.19" />
                    <SPLIT distance="150" swimtime="00:01:37.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:51.39" eventid="1971" heatid="4826" lane="4" />
                <ENTRY entrytime="00:00:56.10" eventid="2013" heatid="4873" lane="3" />
                <ENTRY entrytime="00:00:26.80" eventid="2103" heatid="4946" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Kevin" gender="M" lastname="Kertész" nation="GER" license="391557" athleteid="4188">
              <RESULTS>
                <RESULT eventid="1749" points="441" swimtime="00:02:10.50" resultid="4189" heatid="4677" lane="4" entrytime="00:02:08.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:02.73" />
                    <SPLIT distance="150" swimtime="00:01:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="417" swimtime="00:02:26.71" resultid="4190" heatid="4750" lane="6" entrytime="00:02:25.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:53.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:00.17" eventid="1971" heatid="4813" lane="6" />
                <ENTRY entrytime="00:04:39.87" eventid="2075" heatid="4906" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Hanna" gender="F" lastname="Krauß" nation="GER" license="145397" athleteid="4193">
              <RESULTS>
                <RESULT eventid="1771" points="570" swimtime="00:05:12.85" resultid="4194" heatid="4708" lane="5" entrytime="00:05:09.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                    <SPLIT distance="150" swimtime="00:01:49.20" />
                    <SPLIT distance="200" swimtime="00:02:29.51" />
                    <SPLIT distance="250" swimtime="00:03:15.24" />
                    <SPLIT distance="300" swimtime="00:04:01.47" />
                    <SPLIT distance="350" swimtime="00:04:37.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="652" swimtime="00:04:30.33" resultid="4195" heatid="4763" lane="2" entrytime="00:04:35.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                    <SPLIT distance="100" swimtime="00:01:05.35" />
                    <SPLIT distance="150" swimtime="00:01:39.54" />
                    <SPLIT distance="200" swimtime="00:02:13.82" />
                    <SPLIT distance="250" swimtime="00:02:47.87" />
                    <SPLIT distance="300" swimtime="00:03:22.48" />
                    <SPLIT distance="350" swimtime="00:03:56.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="480" swimtime="00:00:31.13" resultid="4196" heatid="4798" lane="6" entrytime="00:00:30.97" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.16" eventid="1978" heatid="4838" lane="1" />
                <ENTRY entrytime="00:09:29.29" eventid="2020" heatid="4876" lane="6">
                  <MEETINFO qualificationtime="00:09:29.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Katrin" gender="F" lastname="Krauß" nation="GER" license="162021" athleteid="4199">
              <RESULTS>
                <RESULT eventid="1059" points="527" swimtime="00:01:03.02" resultid="4200" heatid="4673" lane="5" entrytime="00:00:59.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="569" swimtime="00:04:42.85" resultid="4201" heatid="4762" lane="2" entrytime="00:04:40.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:39.28" />
                    <SPLIT distance="200" swimtime="00:02:15.37" />
                    <SPLIT distance="250" swimtime="00:02:52.34" />
                    <SPLIT distance="300" swimtime="00:03:29.79" />
                    <SPLIT distance="350" swimtime="00:04:06.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.67" eventid="1978" heatid="4836" lane="1" />
                <ENTRY entrytime="00:00:27.84" eventid="2082" heatid="4922" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Dorothea" gender="F" lastname="Rupprecht" nation="GER" license="271055" athleteid="4205">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.36" eventid="2082" heatid="4915" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia-Sophia" gender="F" lastname="Scheuermann" nation="GER" license="187882" athleteid="4209">
              <RESULTS>
                <RESULT eventid="1771" points="483" swimtime="00:05:30.58" resultid="4210" heatid="4706" lane="1" entrytime="00:05:34.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:17.55" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                    <SPLIT distance="200" swimtime="00:02:43.46" />
                    <SPLIT distance="250" swimtime="00:03:30.59" />
                    <SPLIT distance="300" swimtime="00:04:17.90" />
                    <SPLIT distance="350" swimtime="00:04:54.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Bastian" gender="M" lastname="Schorr" nation="GER" license="137664" athleteid="4212">
              <RESULTS>
                <RESULT eventid="1749" points="615" swimtime="00:01:56.80" resultid="4213" heatid="4684" lane="3" entrytime="00:01:50.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                    <SPLIT distance="100" swimtime="00:00:56.54" />
                    <SPLIT distance="150" swimtime="00:01:26.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="549" swimtime="00:00:59.14" resultid="4214" heatid="4715" lane="3" entrytime="00:00:56.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="556" swimtime="00:00:24.63" resultid="4215" heatid="4776" lane="2" entrytime="00:00:23.65" />
                <RESULT eventid="5369" points="564" swimtime="00:00:58.61" resultid="5377" heatid="5378" lane="4" entrytime="00:00:59.14" />
                <RESULT eventid="1898" points="548" swimtime="00:00:59.16" resultid="5464" heatid="5465" lane="6" entrytime="00:00:59.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:51.17" eventid="1971" heatid="4827" lane="4" />
                <ENTRY entrytime="00:00:58.85" eventid="2027" heatid="4879" lane="3" />
                <ENTRY entrytime="00:00:25.49" eventid="2103" heatid="4945" lane="3" />
                <ENTRY entrytime="00:01:56.80" eventid="1870" heatid="5342" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Corina" gender="F" lastname="Schwandner" nation="GER" license="233736" athleteid="4219">
              <RESULTS>
                <RESULT eventid="1059" points="486" swimtime="00:01:04.73" resultid="4220" heatid="4665" lane="5" entrytime="00:01:03.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:19.38" eventid="1978" heatid="4831" lane="2" />
                <ENTRY entrytime="00:00:28.96" eventid="2082" heatid="4917" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Martin" gender="M" lastname="Spörlein" nation="GER" license="169787" athleteid="4223">
              <RESULTS>
                <RESULT eventid="1834" points="603" swimtime="00:00:23.97" resultid="4224" heatid="4776" lane="4" entrytime="00:00:23.36" />
                <RESULT eventid="1947" points="616" swimtime="00:00:23.81" resultid="5472" heatid="5478" lane="3" entrytime="00:00:23.97" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.66" eventid="1971" heatid="4823" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Fabienne" gender="F" lastname="Wenske" nation="GER" license="287819" swrid="5195433" athleteid="4226">
              <RESULTS>
                <RESULT eventid="1059" points="467" swimtime="00:01:05.58" resultid="4227" heatid="4664" lane="1" entrytime="00:01:04.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1771" points="471" swimtime="00:05:33.44" resultid="4228" heatid="4705" lane="4" entrytime="00:05:39.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:02:01.57" />
                    <SPLIT distance="200" swimtime="00:02:44.15" />
                    <SPLIT distance="250" swimtime="00:03:31.46" />
                    <SPLIT distance="300" swimtime="00:04:21.45" />
                    <SPLIT distance="350" swimtime="00:04:58.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="566" swimtime="00:04:43.45" resultid="4229" heatid="4761" lane="4" entrytime="00:04:45.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:43.51" />
                    <SPLIT distance="200" swimtime="00:02:19.78" />
                    <SPLIT distance="250" swimtime="00:02:55.90" />
                    <SPLIT distance="300" swimtime="00:03:32.10" />
                    <SPLIT distance="350" swimtime="00:04:08.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="569" swimtime="00:18:29.28" resultid="4230" heatid="4803" lane="1" entrytime="00:18:55.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                    <SPLIT distance="150" swimtime="00:01:46.92" />
                    <SPLIT distance="200" swimtime="00:02:23.90" />
                    <SPLIT distance="250" swimtime="00:03:00.98" />
                    <SPLIT distance="300" swimtime="00:03:38.04" />
                    <SPLIT distance="350" swimtime="00:04:15.25" />
                    <SPLIT distance="400" swimtime="00:04:52.55" />
                    <SPLIT distance="450" swimtime="00:05:29.75" />
                    <SPLIT distance="500" swimtime="00:06:06.84" />
                    <SPLIT distance="550" swimtime="00:06:44.28" />
                    <SPLIT distance="600" swimtime="00:07:21.58" />
                    <SPLIT distance="650" swimtime="00:07:58.98" />
                    <SPLIT distance="700" swimtime="00:08:36.12" />
                    <SPLIT distance="750" swimtime="00:09:13.50" />
                    <SPLIT distance="800" swimtime="00:09:50.72" />
                    <SPLIT distance="850" swimtime="00:10:28.02" />
                    <SPLIT distance="900" swimtime="00:11:05.23" />
                    <SPLIT distance="950" swimtime="00:11:42.73" />
                    <SPLIT distance="1000" swimtime="00:12:19.84" />
                    <SPLIT distance="1050" swimtime="00:12:56.90" />
                    <SPLIT distance="1100" swimtime="00:13:34.14" />
                    <SPLIT distance="1150" swimtime="00:14:11.61" />
                    <SPLIT distance="1200" swimtime="00:14:48.84" />
                    <SPLIT distance="1250" swimtime="00:15:26.04" />
                    <SPLIT distance="1300" swimtime="00:16:03.25" />
                    <SPLIT distance="1350" swimtime="00:16:40.19" />
                    <SPLIT distance="1400" swimtime="00:17:17.17" />
                    <SPLIT distance="1450" swimtime="00:17:53.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:16.87" eventid="1978" heatid="4832" lane="2" />
                <ENTRY entrytime="00:02:36.18" eventid="2055" heatid="4899" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Simon" gender="M" lastname="Wicht" nation="GER" license="233738" athleteid="4233">
              <RESULTS>
                <RESULT eventid="1778" points="553" swimtime="00:00:58.98" resultid="4234" heatid="4714" lane="4" entrytime="00:00:57.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="517" swimtime="00:00:27.68" resultid="4235" heatid="4742" lane="4" entrytime="00:00:27.43" />
                <RESULT eventid="1848" points="537" swimtime="00:02:09.92" resultid="4236" heatid="4789" lane="3" entrytime="00:02:07.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:03.53" />
                    <SPLIT distance="150" swimtime="00:01:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2013" status="WDR" swimtime="00:00:00.00" resultid="4237" heatid="4873" lane="4" entrytime="00:00:58.80" />
                <RESULT eventid="2041" status="WDR" swimtime="00:00:00.00" resultid="4238" heatid="4893" lane="4" entrytime="00:02:09.16" />
                <RESULT eventid="2103" status="WDR" swimtime="00:00:00.00" resultid="4239" heatid="4947" lane="1" entrytime="00:00:26.59" />
                <RESULT eventid="1912" points="519" swimtime="00:00:27.64" resultid="5410" heatid="4744" lane="6" entrytime="00:00:27.68" />
                <RESULT eventid="1898" points="562" swimtime="00:00:58.68" resultid="5462" heatid="5465" lane="5" entrytime="00:00:58.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="541" swimtime="00:02:09.63" resultid="5494" heatid="4792" lane="2" entrytime="00:02:09.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="150" swimtime="00:01:36.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="580" swimtime="00:01:48.49" resultid="4240" heatid="4806" lane="5" entrytime="00:01:46.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="100" swimtime="00:00:59.27" />
                    <SPLIT distance="150" swimtime="00:01:25.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4181" number="1" />
                    <RELAYPOSITION athleteid="4233" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="4212" number="3" reactiontime="+33" />
                    <RELAYPOSITION athleteid="4223" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:36.30" eventid="2232" heatid="4812" lane="5" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5095" nation="GER" region="02" clubid="2755" name="SG Frankenhöhe">
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Johannes" gender="M" lastname="Heinz" nation="GER" license="311886" athleteid="2756">
              <RESULTS>
                <RESULT eventid="1763" points="565" swimtime="00:01:07.26" resultid="2757" heatid="4700" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.99" eventid="1985" heatid="4845" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5715" nation="GER" region="02" clubid="3423" name="SG Gundelfingen">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-01" firstname="Charlotte" gender="F" lastname="Joas" nation="GER" license="208201" athleteid="3424">
              <RESULTS>
                <RESULT eventid="1756" points="522" swimtime="00:00:35.75" resultid="3425" heatid="4690" lane="2" entrytime="00:00:36.19" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:19.36" eventid="1992" heatid="4852" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Franziska" gender="F" lastname="Joas" nation="GER" license="155298" athleteid="3427">
              <RESULTS>
                <RESULT eventid="1059" points="525" swimtime="00:01:03.10" resultid="3428" heatid="4667" lane="2" entrytime="00:01:02.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="543" swimtime="00:00:35.28" resultid="3429" heatid="4693" lane="6" entrytime="00:00:35.26" />
                <RESULT eventid="1799" points="512" swimtime="00:01:10.80" resultid="3430" heatid="4731" lane="1" entrytime="00:01:12.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="482" swimtime="00:00:31.09" resultid="3431" heatid="4798" lane="4" entrytime="00:00:30.74" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:18.02" eventid="1992" heatid="4853" lane="3" />
                <ENTRY entrytime="00:00:28.53" eventid="2082" heatid="4919" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5068" nation="GER" region="02" clubid="2406" name="SG Haßberge">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Jonathan" gender="M" lastname="Bischoff" nation="GER" license="260458" athleteid="2407">
              <RESULTS>
                <RESULT eventid="1763" points="455" swimtime="00:01:12.25" resultid="2408" heatid="4697" lane="4" entrytime="00:01:12.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="447" swimtime="00:00:26.48" resultid="2409" heatid="4767" lane="3" entrytime="00:00:26.59" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.35" eventid="1985" heatid="4843" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6768" nation="GER" region="02" clubid="3796" name="SG Mittelfranken">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Varinka" gender="F" lastname="Albert" nation="GER" license="210745" swrid="4193873" athleteid="3801">
              <RESULTS>
                <RESULT eventid="1785" points="578" swimtime="00:01:06.06" resultid="3802" heatid="4723" lane="4" entrytime="00:01:04.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="531" swimtime="00:00:30.10" resultid="3803" heatid="4961" lane="4" entrytime="00:00:28.41" />
                <RESULT eventid="1891" points="591" swimtime="00:01:05.57" resultid="5385" heatid="5391" lane="3" entrytime="00:01:06.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="555" swimtime="00:00:29.66" resultid="5515" heatid="5517" lane="1" entrytime="00:00:30.10" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:04.14" eventid="2006" heatid="4865" lane="4" />
                <ENTRY entrytime="00:00:29.18" eventid="2034" heatid="4889" lane="3" />
                <ENTRY entrytime="00:00:28.13" eventid="2082" heatid="4923" lane="6" />
                <ENTRY entrytime="00:02:18.88" eventid="2096" heatid="4937" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Cindy" gender="F" lastname="Blum" nation="GER" license="291192" athleteid="3808">
              <RESULTS>
                <RESULT eventid="1059" points="552" swimtime="00:01:02.05" resultid="3809" heatid="4671" lane="6" entrytime="00:01:01.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="445" swimtime="00:01:12.04" resultid="3810" heatid="4719" lane="5" entrytime="00:01:12.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="531" swimtime="00:04:49.61" resultid="3811" heatid="4761" lane="2" entrytime="00:04:46.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:06.35" />
                    <SPLIT distance="150" swimtime="00:01:43.25" />
                    <SPLIT distance="200" swimtime="00:02:20.70" />
                    <SPLIT distance="250" swimtime="00:02:57.94" />
                    <SPLIT distance="300" swimtime="00:03:35.65" />
                    <SPLIT distance="350" swimtime="00:04:13.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:14.65" eventid="1978" heatid="4834" lane="1" />
                <ENTRY entrytime="00:10:02.72" eventid="2020" heatid="4875" lane="6">
                  <MEETINFO qualificationtime="00:10:02.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.04" eventid="2082" heatid="4922" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Bruno" gender="M" lastname="Budde" nation="GER" license="272165" athleteid="3816">
              <RESULTS>
                <RESULT eventid="1749" points="477" swimtime="00:02:07.15" resultid="3817" heatid="4679" lane="6" entrytime="00:02:05.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="100" swimtime="00:01:00.71" />
                    <SPLIT distance="150" swimtime="00:01:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1792" points="512" swimtime="00:17:40.02" resultid="3818" heatid="4726" lane="4" entrytime="00:17:44.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:03.22" />
                    <SPLIT distance="150" swimtime="00:01:37.29" />
                    <SPLIT distance="200" swimtime="00:02:11.31" />
                    <SPLIT distance="250" swimtime="00:02:45.53" />
                    <SPLIT distance="300" swimtime="00:03:20.39" />
                    <SPLIT distance="350" swimtime="00:03:55.46" />
                    <SPLIT distance="400" swimtime="00:04:30.75" />
                    <SPLIT distance="450" swimtime="00:05:05.51" />
                    <SPLIT distance="500" swimtime="00:05:40.69" />
                    <SPLIT distance="550" swimtime="00:06:16.13" />
                    <SPLIT distance="600" swimtime="00:06:52.18" />
                    <SPLIT distance="650" swimtime="00:07:28.59" />
                    <SPLIT distance="700" swimtime="00:08:04.50" />
                    <SPLIT distance="750" swimtime="00:08:41.12" />
                    <SPLIT distance="800" swimtime="00:09:17.87" />
                    <SPLIT distance="850" swimtime="00:09:54.10" />
                    <SPLIT distance="900" swimtime="00:10:30.16" />
                    <SPLIT distance="950" swimtime="00:11:05.69" />
                    <SPLIT distance="1000" swimtime="00:11:41.98" />
                    <SPLIT distance="1050" swimtime="00:12:18.71" />
                    <SPLIT distance="1100" swimtime="00:12:55.30" />
                    <SPLIT distance="1150" swimtime="00:13:31.70" />
                    <SPLIT distance="1200" swimtime="00:14:07.77" />
                    <SPLIT distance="1250" swimtime="00:14:43.81" />
                    <SPLIT distance="1300" swimtime="00:15:19.89" />
                    <SPLIT distance="1350" swimtime="00:15:55.16" />
                    <SPLIT distance="1400" swimtime="00:16:31.43" />
                    <SPLIT distance="1450" swimtime="00:17:06.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="411" swimtime="00:02:27.35" resultid="3819" heatid="4752" lane="2" entrytime="00:02:19.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                    <SPLIT distance="150" swimtime="00:01:54.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:57.75" eventid="1999" heatid="4861" lane="6" />
                <ENTRY entrytime="00:02:19.25" eventid="2041" heatid="4891" lane="3" />
                <ENTRY entrytime="00:00:27.86" eventid="2103" heatid="4942" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Leon" gender="M" lastname="Dresel" nation="GER" license="260105" athleteid="3823">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.09" eventid="1971" heatid="4813" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Justin-Joy" gender="M" lastname="Dutschke" nation="GER" license="293147" athleteid="3825">
              <RESULTS>
                <RESULT eventid="1763" points="569" swimtime="00:01:07.09" resultid="3826" heatid="4699" lane="2" entrytime="00:01:10.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="453" swimtime="00:02:22.71" resultid="3827" heatid="4749" lane="3" entrytime="00:02:26.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="100" swimtime="00:01:09.91" />
                    <SPLIT distance="150" swimtime="00:01:49.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.93" eventid="1971" heatid="4816" lane="2" />
                <ENTRY entrytime="00:00:32.51" eventid="1985" heatid="4843" lane="5" />
                <ENTRY entrytime="00:02:34.03" eventid="2089" heatid="4927" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Dominique" gender="F" lastname="Freisleben" nation="GER" license="242096" athleteid="3835">
              <RESULTS>
                <RESULT eventid="1059" points="554" swimtime="00:01:01.95" resultid="3836" heatid="4671" lane="1" entrytime="00:01:01.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="571" swimtime="00:04:42.67" resultid="3837" heatid="4763" lane="5" entrytime="00:04:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="150" swimtime="00:01:40.08" />
                    <SPLIT distance="200" swimtime="00:02:15.59" />
                    <SPLIT distance="250" swimtime="00:02:52.03" />
                    <SPLIT distance="300" swimtime="00:03:28.86" />
                    <SPLIT distance="350" swimtime="00:04:06.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="580" swimtime="00:18:22.37" resultid="3838" heatid="4803" lane="3" entrytime="00:18:26.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:43.14" />
                    <SPLIT distance="200" swimtime="00:02:18.92" />
                    <SPLIT distance="250" swimtime="00:02:55.19" />
                    <SPLIT distance="300" swimtime="00:03:31.61" />
                    <SPLIT distance="350" swimtime="00:04:08.02" />
                    <SPLIT distance="400" swimtime="00:04:44.73" />
                    <SPLIT distance="450" swimtime="00:05:21.69" />
                    <SPLIT distance="500" swimtime="00:05:58.58" />
                    <SPLIT distance="550" swimtime="00:06:35.84" />
                    <SPLIT distance="600" swimtime="00:07:13.12" />
                    <SPLIT distance="650" swimtime="00:07:50.34" />
                    <SPLIT distance="700" swimtime="00:08:27.74" />
                    <SPLIT distance="750" swimtime="00:09:04.58" />
                    <SPLIT distance="800" swimtime="00:09:41.80" />
                    <SPLIT distance="850" swimtime="00:10:18.90" />
                    <SPLIT distance="900" swimtime="00:10:56.10" />
                    <SPLIT distance="950" swimtime="00:11:33.49" />
                    <SPLIT distance="1000" swimtime="00:12:10.77" />
                    <SPLIT distance="1050" swimtime="00:12:48.51" />
                    <SPLIT distance="1100" swimtime="00:13:25.85" />
                    <SPLIT distance="1150" swimtime="00:14:03.17" />
                    <SPLIT distance="1200" swimtime="00:14:40.43" />
                    <SPLIT distance="1250" swimtime="00:15:17.83" />
                    <SPLIT distance="1300" swimtime="00:15:55.07" />
                    <SPLIT distance="1350" swimtime="00:16:32.38" />
                    <SPLIT distance="1400" swimtime="00:17:09.68" />
                    <SPLIT distance="1450" swimtime="00:17:46.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:12.00" eventid="1978" heatid="4835" lane="3" />
                <ENTRY entrytime="00:09:30.00" eventid="2020" heatid="4875" lane="3">
                  <MEETINFO qualificationtime="00:09:30.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.00" eventid="2082" heatid="4921" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Mareike" gender="F" lastname="Förster" nation="GER" license="183768" athleteid="3831">
              <RESULTS>
                <RESULT eventid="1756" points="599" swimtime="00:00:34.16" resultid="3832" heatid="4694" lane="4" entrytime="00:00:33.22" />
                <RESULT eventid="1799" points="621" swimtime="00:01:06.41" resultid="3833" heatid="4735" lane="4" entrytime="00:01:06.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="624" swimtime="00:02:37.44" resultid="3834" heatid="4783" lane="3" entrytime="00:02:28.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:16.10" />
                    <SPLIT distance="150" swimtime="00:01:55.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1877" points="577" swimtime="00:00:34.58" resultid="5350" heatid="5355" lane="4" entrytime="00:00:34.16" />
                <RESULT eventid="1919" points="618" swimtime="00:01:06.53" resultid="5394" heatid="4737" lane="2" entrytime="00:01:06.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1954" points="607" swimtime="00:02:38.93" resultid="5481" heatid="4785" lane="2" entrytime="00:02:37.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Selina" gender="F" lastname="Herzog" nation="GER" license="274715" athleteid="3842">
              <RESULTS>
                <RESULT eventid="1756" points="434" swimtime="00:00:38.02" resultid="3843" heatid="4688" lane="4" entrytime="00:00:37.18" />
                <RESULT eventid="1841" points="425" swimtime="00:02:58.87" resultid="3844" heatid="4779" lane="4" entrytime="00:02:57.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:25.05" />
                    <SPLIT distance="150" swimtime="00:02:12.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="393" swimtime="00:00:33.26" resultid="3845" heatid="4794" lane="2" entrytime="00:00:32.03" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:22.51" eventid="1992" heatid="4850" lane="5" />
                <ENTRY entrytime="00:01:10.47" eventid="2006" heatid="4864" lane="6" />
                <ENTRY entrytime="00:02:39.35" eventid="2055" heatid="4896" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Benno" gender="M" lastname="Hingler" nation="GER" license="242439" athleteid="3849">
              <RESULTS>
                <RESULT eventid="1763" points="480" swimtime="00:01:11.01" resultid="3850" heatid="4698" lane="2" entrytime="00:01:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="421" swimtime="00:00:29.63" resultid="3851" heatid="4740" lane="1" entrytime="00:00:29.84" />
                <RESULT eventid="1820" points="452" swimtime="00:02:22.75" resultid="3852" heatid="4751" lane="2" entrytime="00:02:22.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                    <SPLIT distance="100" swimtime="00:01:07.33" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="494" swimtime="00:00:25.62" resultid="3853" heatid="4769" lane="4" entrytime="00:00:26.11" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.72" eventid="1985" heatid="4844" lane="2" />
                <ENTRY entrytime="00:01:03.02" eventid="2027" heatid="4881" lane="1" />
                <ENTRY entrytime="00:02:37.57" eventid="2089" heatid="4926" lane="2" />
                <ENTRY entrytime="00:00:27.36" eventid="2103" heatid="4944" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Hannah" gender="F" lastname="Hofmockel" nation="GER" license="256656" athleteid="3858">
              <RESULTS>
                <RESULT eventid="1756" points="535" swimtime="00:00:35.47" resultid="3859" heatid="4694" lane="5" entrytime="00:00:34.10" />
                <RESULT eventid="1799" points="542" swimtime="00:01:09.48" resultid="3860" heatid="4734" lane="2" entrytime="00:01:08.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="525" swimtime="00:02:46.79" resultid="3861" heatid="4783" lane="4" entrytime="00:02:39.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:19.98" />
                    <SPLIT distance="150" swimtime="00:02:03.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1919" points="547" swimtime="00:01:09.26" resultid="5397" heatid="4737" lane="6" entrytime="00:01:09.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:14.65" eventid="1992" heatid="4855" lane="4" />
                <ENTRY entrytime="NT" eventid="2020" status="RJC" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Simon" gender="M" lastname="Jonscher" nation="GER" license="271097" athleteid="3865">
              <RESULTS>
                <RESULT eventid="1749" points="540" swimtime="00:02:01.98" resultid="3866" heatid="4682" lane="1" entrytime="00:02:00.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="100" swimtime="00:00:58.94" />
                    <SPLIT distance="150" swimtime="00:01:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="465" swimtime="00:01:02.49" resultid="3867" heatid="4712" lane="1" entrytime="00:01:01.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="481" swimtime="00:00:25.85" resultid="3868" heatid="4770" lane="1" entrytime="00:00:26.00" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.47" eventid="1971" heatid="4822" lane="6" />
                <ENTRY entrytime="00:01:04.54" eventid="2013" heatid="4870" lane="6" />
                <ENTRY entrytime="00:00:28.23" eventid="2103" heatid="4941" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Jens" gender="M" lastname="Jüttner" nation="GER" license="179877" athleteid="3872">
              <RESULTS>
                <RESULT eventid="1834" points="525" swimtime="00:00:25.11" resultid="3873" heatid="4771" lane="3" entrytime="00:00:25.59" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Daniela" gender="F" lastname="Karst" nation="GER" license="156320" athleteid="3874">
              <RESULTS>
                <RESULT eventid="1756" status="DNS" swimtime="00:00:00.00" resultid="3875" heatid="4692" lane="3" entrytime="00:00:33.11" />
                <RESULT eventid="1799" status="DNS" swimtime="00:00:00.00" resultid="3876" heatid="4736" lane="4" entrytime="00:01:06.41" />
                <RESULT eventid="1813" status="DNS" swimtime="00:00:00.00" resultid="3877" heatid="4746" lane="3" entrytime="00:02:17.97" />
                <RESULT eventid="1855" status="DNS" swimtime="00:00:00.00" resultid="3878" heatid="4801" lane="4" entrytime="00:00:28.42" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:11.57" eventid="1992" heatid="4857" lane="3" />
                <ENTRY entrytime="00:01:03.15" eventid="2006" heatid="4866" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Kai" gender="M" lastname="Kisberi" nation="GER" license="196491" athleteid="3881">
              <RESULTS>
                <RESULT eventid="1749" points="496" swimtime="00:02:05.45" resultid="3882" heatid="4681" lane="3" entrytime="00:02:01.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                    <SPLIT distance="100" swimtime="00:01:00.08" />
                    <SPLIT distance="150" swimtime="00:01:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="458" swimtime="00:00:26.27" resultid="3883" heatid="4769" lane="2" entrytime="00:00:26.15" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.74" eventid="1971" heatid="4819" lane="2" />
                <ENTRY entrytime="00:04:20.97" eventid="2075" heatid="4909" lane="3" />
                <ENTRY entrytime="NT" eventid="2168" status="RJC" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Daniel" gender="M" lastname="Knorr" nation="GER" license="270253" athleteid="3887">
              <RESULTS>
                <RESULT eventid="1778" points="463" swimtime="00:01:02.61" resultid="3888" heatid="4710" lane="5" entrytime="00:01:03.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="479" swimtime="00:02:20.09" resultid="3889" heatid="4752" lane="6" entrytime="00:02:21.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:03.87" />
                    <SPLIT distance="150" swimtime="00:01:46.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="438" swimtime="00:02:19.08" resultid="3890" heatid="4791" lane="6" entrytime="00:02:15.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:43.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.61" eventid="1971" heatid="4817" lane="1" />
                <ENTRY entrytime="00:01:03.50" eventid="2013" heatid="4870" lane="4" />
                <ENTRY entrytime="00:02:16.82" eventid="2041" heatid="4892" lane="1" />
                <ENTRY entrytime="00:00:28.92" eventid="2103" heatid="4940" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Arthur" gender="M" lastname="Kraft" nation="GER" license="260249" athleteid="3895">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.79" eventid="1971" heatid="4816" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Oliver" gender="M" lastname="Kreißel" nation="GER" license="313677" athleteid="3897">
              <RESULTS>
                <RESULT eventid="1763" points="372" swimtime="00:01:17.29" resultid="3898" heatid="4696" lane="2" entrytime="00:01:14.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:33.20" eventid="1985" heatid="4842" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Denis" gender="M" lastname="Kremer" nation="GER" license="302575" athleteid="3900">
              <RESULTS>
                <RESULT eventid="1778" points="496" swimtime="00:01:01.18" resultid="3901" heatid="4709" lane="2" entrytime="00:01:04.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="462" swimtime="00:00:28.73" resultid="3902" heatid="4743" lane="6" entrytime="00:00:29.10" />
                <RESULT eventid="1834" points="491" swimtime="00:00:25.67" resultid="3903" heatid="4768" lane="3" entrytime="00:00:26.33" />
                <RESULT eventid="1848" points="412" swimtime="00:02:21.90" resultid="3904" heatid="4788" lane="1" entrytime="00:02:19.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:59.48" eventid="1971" heatid="4814" lane="2" />
                <ENTRY entrytime="00:01:04.05" eventid="2013" heatid="4870" lane="5" />
                <ENTRY entrytime="00:01:05.93" eventid="2027" heatid="4877" lane="3" />
                <ENTRY entrytime="00:00:27.03" eventid="2103" heatid="4945" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Elija" gender="M" lastname="Krewer" nation="GER" license="253067" athleteid="3909">
              <ENTRIES>
                <ENTRY entrytime="00:04:36.49" eventid="2075" heatid="4907" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Liv" gender="F" lastname="Krumme" nation="GER" license="281732" athleteid="3911">
              <RESULTS>
                <RESULT eventid="1059" points="537" swimtime="00:01:02.60" resultid="3912" heatid="4670" lane="4" entrytime="00:01:01.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="473" swimtime="00:01:10.60" resultid="3913" heatid="4721" lane="4" entrytime="00:01:08.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:15.44" eventid="1978" heatid="4833" lane="2" />
                <ENTRY entrytime="00:00:32.77" eventid="2034" heatid="4886" lane="5" />
                <ENTRY entrytime="00:02:35.02" eventid="2055" heatid="4900" lane="2" />
                <ENTRY entrytime="00:00:28.93" eventid="2082" heatid="4917" lane="3" />
                <ENTRY entrytime="00:02:25.59" eventid="2096" heatid="4935" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Kellie" gender="F" lastname="Messel" nation="GER" license="321746" athleteid="3919">
              <RESULTS>
                <RESULT eventid="1059" points="475" swimtime="00:01:05.23" resultid="3920" heatid="4665" lane="6" entrytime="00:01:03.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="444" swimtime="00:00:37.73" resultid="3921" heatid="4687" lane="6" entrytime="00:00:38.03" />
                <RESULT eventid="1827" points="545" swimtime="00:04:47.07" resultid="3922" heatid="4759" lane="4" entrytime="00:04:54.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:45.27" />
                    <SPLIT distance="200" swimtime="00:02:22.04" />
                    <SPLIT distance="250" swimtime="00:02:58.32" />
                    <SPLIT distance="300" swimtime="00:03:35.34" />
                    <SPLIT distance="350" swimtime="00:04:12.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="482" swimtime="00:02:51.63" resultid="3923" heatid="4780" lane="5" entrytime="00:02:53.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:23.32" />
                    <SPLIT distance="150" swimtime="00:02:07.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:20.61" eventid="1992" heatid="4851" lane="1" />
                <ENTRY entrytime="00:02:40.27" eventid="2055" heatid="4896" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Michelle" gender="F" lastname="Messel" nation="GER" license="196996" athleteid="3926">
              <RESULTS>
                <RESULT eventid="1813" points="587" swimtime="00:02:22.83" resultid="3927" heatid="4745" lane="3" entrytime="00:02:18.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="600" swimtime="00:00:28.89" resultid="3928" heatid="4800" lane="3" entrytime="00:00:28.23" />
                <RESULT eventid="1933" points="598" swimtime="00:02:21.95" resultid="5419" heatid="4748" lane="4" entrytime="00:02:22.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                    <SPLIT distance="150" swimtime="00:01:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="597" swimtime="00:00:28.95" resultid="5507" heatid="4802" lane="2" entrytime="00:00:28.89" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:03.50" eventid="2006" heatid="4865" lane="3" />
                <ENTRY entrytime="00:00:31.80" eventid="2034" heatid="4887" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Christoph" gender="M" lastname="Mooser" nation="GER" license="240870" athleteid="3931">
              <RESULTS>
                <RESULT eventid="1763" points="580" swimtime="00:01:06.66" resultid="3932" heatid="4701" lane="1" entrytime="00:01:06.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="488" swimtime="00:00:28.22" resultid="3933" heatid="4741" lane="2" entrytime="00:00:28.05" />
                <RESULT eventid="1820" points="551" swimtime="00:02:13.66" resultid="3934" heatid="4756" lane="1" entrytime="00:02:11.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:04.72" />
                    <SPLIT distance="150" swimtime="00:01:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="481" swimtime="00:02:14.80" resultid="3935" heatid="4789" lane="5" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.31" />
                    <SPLIT distance="100" swimtime="00:01:05.96" />
                    <SPLIT distance="150" swimtime="00:01:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1912" points="492" swimtime="00:00:28.13" resultid="5415" heatid="5417" lane="1" entrytime="00:00:28.22" />
                <RESULT eventid="1961" points="512" swimtime="00:02:12.03" resultid="5498" heatid="5504" lane="3" entrytime="00:02:14.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="150" swimtime="00:01:38.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.09" eventid="1985" heatid="4848" lane="1" />
                <ENTRY entrytime="00:01:00.21" eventid="2013" heatid="4871" lane="4" />
                <ENTRY entrytime="00:02:23.26" eventid="2089" heatid="4929" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Jonas" gender="M" lastname="Mursak" nation="GER" license="196445" athleteid="3939">
              <RESULTS>
                <RESULT eventid="1763" points="622" swimtime="00:01:05.14" resultid="3940" heatid="4703" lane="1" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="518" swimtime="00:02:16.48" resultid="3941" heatid="4754" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:44.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1884" points="626" swimtime="00:01:04.99" resultid="5366" heatid="5368" lane="1" entrytime="00:01:05.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.43" eventid="1985" heatid="4848" lane="6" />
                <ENTRY entrytime="00:00:59.94" eventid="2027" heatid="4881" lane="2" />
                <ENTRY entrytime="00:02:22.50" eventid="2089" heatid="4930" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lisa" gender="F" lastname="Mursak" nation="GER" license="196457" athleteid="3945">
              <RESULTS>
                <RESULT eventid="1785" points="614" swimtime="00:01:04.72" resultid="3946" heatid="4723" lane="3" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="511" swimtime="00:00:30.48" resultid="3947" heatid="4797" lane="2" entrytime="00:00:31.03" />
                <RESULT eventid="1891" points="623" swimtime="00:01:04.42" resultid="5381" heatid="4725" lane="2" entrytime="00:01:04.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.90" eventid="2034" heatid="4888" lane="3" />
                <ENTRY entrytime="00:02:18.00" eventid="2096" heatid="4935" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Katja" gender="F" lastname="Neousypin" nation="GER" license="281139" athleteid="3950">
              <RESULTS>
                <RESULT eventid="1756" points="552" swimtime="00:00:35.10" resultid="3951" heatid="4694" lane="1" entrytime="00:00:34.63" />
                <RESULT eventid="1771" points="469" swimtime="00:05:33.76" resultid="3952" heatid="4706" lane="5" entrytime="00:05:34.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                    <SPLIT distance="150" swimtime="00:02:01.92" />
                    <SPLIT distance="200" swimtime="00:02:44.71" />
                    <SPLIT distance="250" swimtime="00:03:30.88" />
                    <SPLIT distance="300" swimtime="00:04:18.45" />
                    <SPLIT distance="350" swimtime="00:04:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="509" swimtime="00:02:48.48" resultid="3953" heatid="4784" lane="5" entrytime="00:02:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:02:05.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="445" swimtime="00:00:31.91" resultid="3954" heatid="4796" lane="2" entrytime="00:00:31.41" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:15.40" eventid="1992" heatid="4857" lane="2" />
                <ENTRY entrytime="00:01:10.46" eventid="2006" heatid="4864" lane="1" />
                <ENTRY entrytime="00:02:33.79" eventid="2055" heatid="4901" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Tanja" gender="F" lastname="Neubert" nation="GER" license="274074" athleteid="3958">
              <RESULTS>
                <RESULT eventid="1756" points="514" swimtime="00:00:35.94" resultid="3959" heatid="4690" lane="1" entrytime="00:00:36.43" />
                <RESULT eventid="1841" points="531" swimtime="00:02:46.10" resultid="3960" heatid="4784" lane="1" entrytime="00:02:45.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:21.07" />
                    <SPLIT distance="150" swimtime="00:02:04.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1954" points="509" swimtime="00:02:48.48" resultid="5490" heatid="5491" lane="6" entrytime="00:02:46.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:20.67" />
                    <SPLIT distance="150" swimtime="00:02:05.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:16.84" eventid="1992" heatid="4856" lane="6" />
                <ENTRY entrytime="00:02:38.75" eventid="2055" heatid="4897" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Daniela" gender="F" lastname="Neubig" nation="GER" license="169855" athleteid="3963">
              <RESULTS>
                <RESULT eventid="1771" points="631" swimtime="00:05:02.37" resultid="3964" heatid="4708" lane="4" entrytime="00:04:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                    <SPLIT distance="150" swimtime="00:01:47.76" />
                    <SPLIT distance="200" swimtime="00:02:24.85" />
                    <SPLIT distance="250" swimtime="00:03:07.72" />
                    <SPLIT distance="300" swimtime="00:03:50.79" />
                    <SPLIT distance="350" swimtime="00:04:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="551" swimtime="00:02:44.11" resultid="3965" heatid="4784" lane="2" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                    <SPLIT distance="100" swimtime="00:01:19.14" />
                    <SPLIT distance="150" swimtime="00:02:01.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1954" points="560" swimtime="00:02:43.24" resultid="5488" heatid="5491" lane="5" entrytime="00:02:44.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:18.54" />
                    <SPLIT distance="150" swimtime="00:02:00.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:15.77" eventid="1992" heatid="4857" lane="5" />
                <ENTRY entrytime="00:02:23.50" eventid="2055" heatid="4904" lane="2" />
                <ENTRY entrytime="00:02:19.50" eventid="2096" heatid="4936" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Jeremias" gender="M" lastname="Pock" nation="GER" license="269306" athleteid="3969">
              <RESULTS>
                <RESULT eventid="1763" points="439" swimtime="00:01:13.14" resultid="3970" heatid="4696" lane="5" entrytime="00:01:14.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="483" swimtime="00:02:19.71" resultid="3971" heatid="4751" lane="6" entrytime="00:02:22.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:47.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="410" swimtime="00:02:22.15" resultid="3972" heatid="4786" lane="3" entrytime="00:02:22.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:45.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:34.35" eventid="1985" heatid="4841" lane="5" />
                <ENTRY entrytime="00:05:05.35" eventid="1999" heatid="4859" lane="3" />
                <ENTRY entrytime="00:02:38.86" eventid="2089" heatid="4926" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Cosima" gender="F" lastname="Rau" nation="GER" license="295229" athleteid="3976">
              <RESULTS>
                <RESULT eventid="1771" points="537" swimtime="00:05:19.21" resultid="3977" heatid="4707" lane="1" entrytime="00:05:27.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:54.96" />
                    <SPLIT distance="200" swimtime="00:02:35.81" />
                    <SPLIT distance="250" swimtime="00:03:19.99" />
                    <SPLIT distance="300" swimtime="00:04:04.42" />
                    <SPLIT distance="350" swimtime="00:04:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="578" swimtime="00:02:41.48" resultid="3978" heatid="4779" lane="1" entrytime="00:03:06.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:02:01.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1954" points="552" swimtime="00:02:43.97" resultid="5485" heatid="5491" lane="3" entrytime="00:02:41.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:18.61" />
                    <SPLIT distance="150" swimtime="00:02:01.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:18.88" eventid="1992" heatid="4853" lane="1" />
                <ENTRY entrytime="00:02:44.43" eventid="2055" heatid="4896" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Andreas" gender="M" lastname="Rein" nation="GER" license="278278" athleteid="3981">
              <RESULTS>
                <RESULT eventid="1749" points="583" swimtime="00:01:58.89" resultid="3982" heatid="4683" lane="5" entrytime="00:01:55.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                    <SPLIT distance="100" swimtime="00:00:57.45" />
                    <SPLIT distance="150" swimtime="00:01:28.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="592" swimtime="00:00:24.12" resultid="3983" heatid="4777" lane="2" entrytime="00:00:23.47" />
                <RESULT eventid="1848" points="499" swimtime="00:02:13.11" resultid="3984" heatid="4790" lane="4" entrytime="00:02:09.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:03.63" />
                    <SPLIT distance="150" swimtime="00:01:38.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1947" points="600" swimtime="00:00:24.02" resultid="5474" heatid="5478" lane="2" entrytime="00:00:24.12" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:51.11" eventid="1971" heatid="4826" lane="3" />
                <ENTRY entrytime="00:01:02.43" eventid="2013" heatid="4872" lane="6" />
                <ENTRY entrytime="00:00:25.54" eventid="2103" heatid="4945" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Ferdinand" gender="M" lastname="Reng" nation="GER" license="188193" athleteid="3988">
              <RESULTS>
                <RESULT eventid="1834" points="631" swimtime="00:00:23.61" resultid="3989" heatid="4777" lane="4" entrytime="00:00:23.25" />
                <RESULT eventid="1947" points="650" swimtime="00:00:23.38" resultid="5469" heatid="4778" lane="5" entrytime="00:00:23.61" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.39" eventid="1971" heatid="4826" lane="1" />
                <ENTRY entrytime="00:00:26.22" eventid="2103" heatid="4947" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Julian" gender="M" lastname="Richter" nation="GER" license="166195" athleteid="3992">
              <RESULTS>
                <RESULT eventid="1778" points="540" swimtime="00:00:59.48" resultid="3993" heatid="4714" lane="2" entrytime="00:00:58.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.84" eventid="2041" heatid="4892" lane="2" />
                <ENTRY entrytime="00:00:27.61" eventid="2103" heatid="4943" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Nikita" gender="M" lastname="Rodenko" nation="GER" license="361022" athleteid="3996">
              <RESULTS>
                <RESULT eventid="1749" points="698" swimtime="00:01:52.00" resultid="3997" heatid="4684" lane="1" entrytime="00:01:56.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="100" swimtime="00:00:55.16" />
                    <SPLIT distance="150" swimtime="00:01:24.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="589" swimtime="00:02:10.76" resultid="3998" heatid="4756" lane="2" entrytime="00:02:08.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                    <SPLIT distance="100" swimtime="00:01:02.43" />
                    <SPLIT distance="150" swimtime="00:01:40.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="619" swimtime="00:02:08.61" resultid="5438" heatid="5442" lane="2" entrytime="00:02:10.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                    <SPLIT distance="100" swimtime="00:01:02.21" />
                    <SPLIT distance="150" swimtime="00:01:38.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:51.15" eventid="1971" heatid="4825" lane="3" />
                <ENTRY entrytime="00:02:12.90" eventid="2041" heatid="4893" lane="5" />
                <ENTRY entrytime="00:08:33.44" eventid="2168" heatid="4809" lane="6">
                  <MEETINFO qualificationtime="00:08:33.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.00" eventid="1870" heatid="4686" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Nele" gender="F" lastname="Rudolph" nation="GER" license="274362" athleteid="4002">
              <RESULTS>
                <RESULT eventid="1059" points="463" swimtime="00:01:05.80" resultid="4003" heatid="4662" lane="4" entrytime="00:01:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Leonie" gender="F" lastname="Sauer" nation="GER" license="289750" athleteid="4004">
              <RESULTS>
                <RESULT eventid="1771" points="451" swimtime="00:05:38.26" resultid="4005" heatid="4706" lane="4" entrytime="00:05:29.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:02:00.05" />
                    <SPLIT distance="200" swimtime="00:02:43.84" />
                    <SPLIT distance="250" swimtime="00:03:31.13" />
                    <SPLIT distance="300" swimtime="00:04:18.98" />
                    <SPLIT distance="350" swimtime="00:04:59.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="439" swimtime="00:02:56.96" resultid="4006" heatid="4779" lane="3" entrytime="00:02:57.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:01:23.90" />
                    <SPLIT distance="150" swimtime="00:02:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="438" swimtime="00:00:32.10" resultid="4007" heatid="4794" lane="3" entrytime="00:00:31.94" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:21.17" eventid="1992" heatid="4851" lane="6" />
                <ENTRY entrytime="00:02:32.69" eventid="2055" heatid="4901" lane="3" />
                <ENTRY entrytime="00:00:30.08" eventid="2082" heatid="4913" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Helene" gender="F" lastname="Schall" nation="GER" license="309209" athleteid="4011">
              <RESULTS>
                <RESULT eventid="1785" points="507" swimtime="00:01:08.98" resultid="4012" heatid="4721" lane="5" entrytime="00:01:09.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="464" swimtime="00:01:13.15" resultid="4013" heatid="4732" lane="2" entrytime="00:01:12.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:20.60" eventid="1978" heatid="4829" lane="3" />
                <ENTRY entrytime="00:00:31.02" eventid="2034" heatid="4889" lane="5" />
                <ENTRY entrytime="00:02:32.04" eventid="2096" heatid="4934" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Ronja" gender="F" lastname="Scharnweber" nation="GER" license="312797" athleteid="4017">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.04" eventid="2082" heatid="4913" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Lars" gender="M" lastname="Schuseil" nation="GER" license="287319" athleteid="4949">
              <RESULTS>
                <RESULT eventid="1749" points="447" swimtime="00:02:09.91" resultid="4950" heatid="4676" lane="3" entrytime="00:02:10.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:03.32" />
                    <SPLIT distance="150" swimtime="00:01:37.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:59.90" eventid="1971" heatid="4813" lane="3" />
                <ENTRY entrytime="00:04:37.87" eventid="2075" heatid="4907" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Alexander" gender="M" lastname="Sinn" nation="GER" license="169871" athleteid="4019">
              <RESULTS>
                <RESULT eventid="1763" points="528" swimtime="00:01:08.77" resultid="4020" heatid="4700" lane="4" entrytime="00:01:07.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="492" swimtime="00:00:25.66" resultid="4021" heatid="4772" lane="6" entrytime="00:00:25.50" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.00" eventid="1985" heatid="4845" lane="4" />
                <ENTRY entrytime="00:02:26.87" eventid="2089" heatid="4930" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Anna Lena" gender="F" lastname="Sinn" nation="GER" license="169870" athleteid="4024">
              <RESULTS>
                <RESULT eventid="1756" points="625" swimtime="00:00:33.67" resultid="4025" heatid="4693" lane="4" entrytime="00:00:33.38" />
                <RESULT eventid="1877" points="611" swimtime="00:00:33.93" resultid="5347" heatid="4695" lane="1" entrytime="00:00:33.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Laura" gender="F" lastname="Steuerl" nation="GER" license="316690" athleteid="4953">
              <RESULTS>
                <RESULT eventid="1059" points="526" swimtime="00:01:03.05" resultid="4954" heatid="4668" lane="2" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1813" points="453" swimtime="00:02:35.72" resultid="4955" heatid="4745" lane="1" entrytime="00:02:39.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:01:55.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="443" swimtime="00:00:31.98" resultid="4956" heatid="4793" lane="2" entrytime="00:00:32.77" />
                <RESULT eventid="1933" points="457" swimtime="00:02:35.28" resultid="5428" heatid="5429" lane="1" entrytime="00:02:35.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:54.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:15.39" eventid="1978" heatid="4833" lane="4" />
                <ENTRY entrytime="NT" eventid="2020" status="RJC" />
                <ENTRY entrytime="00:00:29.28" eventid="2082" heatid="4916" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lorenz" gender="M" lastname="Streicher" nation="GER" license="252860" athleteid="4026">
              <RESULTS>
                <RESULT eventid="1749" points="496" swimtime="00:02:05.53" resultid="4027" heatid="4678" lane="5" entrytime="00:02:06.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="100" swimtime="00:01:00.96" />
                    <SPLIT distance="150" swimtime="00:01:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="444" swimtime="00:01:03.46" resultid="4028" heatid="4709" lane="1" entrytime="00:01:05.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="456" swimtime="00:02:22.43" resultid="4029" heatid="4750" lane="2" entrytime="00:02:24.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:07.25" />
                    <SPLIT distance="150" swimtime="00:01:51.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="422" swimtime="00:02:20.79" resultid="4030" heatid="4787" lane="5" entrytime="00:02:21.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                    <SPLIT distance="150" swimtime="00:01:45.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:05:02.57" eventid="1999" heatid="4860" lane="5" />
                <ENTRY entrytime="00:04:37.27" eventid="2075" heatid="4907" lane="2" />
                <ENTRY entrytime="00:00:29.11" eventid="2103" heatid="4939" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Elena" gender="F" lastname="Tröger" nation="GER" license="307156" athleteid="4034">
              <ENTRIES>
                <ENTRY entrytime="00:02:18.13" eventid="1978" heatid="4832" lane="6" />
                <ENTRY entrytime="00:02:35.10" eventid="2055" heatid="4900" lane="1" />
                <ENTRY entrytime="00:00:29.98" eventid="2082" heatid="4913" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Felicia" gender="F" lastname="Tröger" nation="GER" license="309284" athleteid="4041">
              <RESULTS>
                <RESULT eventid="1756" points="548" swimtime="00:00:35.19" resultid="4042" heatid="4689" lane="4" entrytime="00:00:36.84" />
                <RESULT eventid="1785" points="458" swimtime="00:01:11.36" resultid="4043" heatid="4719" lane="3" entrytime="00:01:11.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="532" swimtime="00:01:09.93" resultid="4044" heatid="4736" lane="6" entrytime="00:01:11.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="486" swimtime="00:02:51.15" resultid="4045" heatid="4780" lane="2" entrytime="00:02:53.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:22.43" />
                    <SPLIT distance="150" swimtime="00:02:08.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="467" swimtime="00:00:31.41" resultid="4046" heatid="4799" lane="6" entrytime="00:00:30.71" />
                <RESULT eventid="1919" points="558" swimtime="00:01:08.82" resultid="5399" heatid="5404" lane="4" entrytime="00:01:09.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:18.79" eventid="1992" heatid="4853" lane="5" />
                <ENTRY entrytime="00:00:34.49" eventid="2034" heatid="4883" lane="2" />
                <ENTRY entrytime="00:02:39.11" eventid="2055" heatid="4897" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Emma" gender="F" lastname="Veit" nation="GER" license="301073" athleteid="4050">
              <RESULTS>
                <RESULT eventid="1059" points="504" swimtime="00:01:03.97" resultid="4051" heatid="4667" lane="6" entrytime="00:01:03.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="464" swimtime="00:01:11.04" resultid="4052" heatid="4720" lane="2" entrytime="00:01:11.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:10.96" eventid="2006" heatid="4863" lane="4" />
                <ENTRY entrytime="00:02:39.17" eventid="2055" heatid="4897" lane="1" />
                <ENTRY entrytime="00:00:29.46" eventid="2082" heatid="4915" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Karla" gender="F" lastname="Völcker" nation="GER" license="216926" athleteid="4056">
              <RESULTS>
                <RESULT eventid="1059" points="558" swimtime="00:01:01.83" resultid="4057" heatid="4669" lane="5" entrytime="00:01:02.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="583" swimtime="00:01:05.86" resultid="4058" heatid="4724" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="500" swimtime="00:00:30.70" resultid="4059" heatid="4798" lane="1" entrytime="00:00:30.93" />
                <RESULT eventid="1891" points="570" swimtime="00:01:06.36" resultid="5383" heatid="4725" lane="1" entrytime="00:01:05.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:15.22" eventid="1978" heatid="4833" lane="3" />
                <ENTRY entrytime="00:00:30.77" eventid="2034" heatid="4887" lane="4" />
                <ENTRY entrytime="00:00:28.48" eventid="2082" heatid="4919" lane="2" />
                <ENTRY entrytime="00:02:21.86" eventid="2096" heatid="4935" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Annalena" gender="F" lastname="Wagner" nation="GER" license="297332" athleteid="4064">
              <RESULTS>
                <RESULT eventid="1059" points="626" swimtime="00:00:59.50" resultid="4065" heatid="4672" lane="2" entrytime="00:00:59.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="623" swimtime="00:01:04.42" resultid="4066" heatid="4722" lane="5" entrytime="00:01:05.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="639" swimtime="00:04:32.25" resultid="4067" heatid="4763" lane="6" entrytime="00:04:39.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                    <SPLIT distance="200" swimtime="00:02:13.88" />
                    <SPLIT distance="250" swimtime="00:02:48.38" />
                    <SPLIT distance="300" swimtime="00:03:23.19" />
                    <SPLIT distance="350" swimtime="00:03:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="633" swimtime="00:00:59.29" resultid="5323" heatid="4675" lane="6" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1891" points="640" swimtime="00:01:03.85" resultid="5380" heatid="4725" lane="4" entrytime="00:01:04.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:13.46" eventid="1978" heatid="4835" lane="6" />
                <ENTRY entrytime="00:00:31.44" eventid="2034" heatid="4887" lane="5" />
                <ENTRY entrytime="00:02:19.84" eventid="2096" heatid="4935" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Rebecca" gender="F" lastname="Walther" nation="GER" license="292203" athleteid="4071">
              <RESULTS>
                <RESULT eventid="1756" points="471" swimtime="00:00:37.00" resultid="4072" heatid="4687" lane="1" entrytime="00:00:37.96" />
                <RESULT eventid="1841" points="445" swimtime="00:02:56.18" resultid="4073" heatid="4779" lane="5" entrytime="00:02:58.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:01:25.36" />
                    <SPLIT distance="150" swimtime="00:02:11.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Deborah" gender="F" lastname="Weber" nation="GER" license="227778" athleteid="4074">
              <RESULTS>
                <RESULT eventid="1813" points="557" swimtime="00:02:25.35" resultid="4075" heatid="4746" lane="2" entrytime="00:02:25.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:48.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="465" swimtime="00:00:31.46" resultid="4076" heatid="4798" lane="5" entrytime="00:00:30.83" />
                <RESULT eventid="1933" points="586" swimtime="00:02:22.88" resultid="5421" heatid="4748" lane="5" entrytime="00:02:25.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:09.03" />
                    <SPLIT distance="150" swimtime="00:01:46.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:07.13" eventid="2006" heatid="4865" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Josefina" gender="F" lastname="Wiesbeck" nation="GER" license="301078" athleteid="4079">
              <RESULTS>
                <RESULT eventid="1813" points="560" swimtime="00:02:25.06" resultid="4080" heatid="4747" lane="5" entrytime="00:02:29.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="477" swimtime="00:00:31.19" resultid="4081" heatid="4795" lane="2" entrytime="00:00:31.67" />
                <RESULT eventid="1933" points="560" swimtime="00:02:25.08" resultid="5420" heatid="4748" lane="2" entrytime="00:02:25.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:08.45" />
                    <SPLIT distance="150" swimtime="00:01:46.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:08.16" eventid="2006" heatid="4866" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="588" swimtime="00:01:48.00" resultid="4083" heatid="4806" lane="2" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                    <SPLIT distance="100" swimtime="00:00:57.27" />
                    <SPLIT distance="150" swimtime="00:01:23.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3931" number="1" />
                    <RELAYPOSITION athleteid="3939" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3996" number="3" reactiontime="+43" />
                    <RELAYPOSITION athleteid="3988" number="4" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:35.00" eventid="2232" heatid="4812" lane="2" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="2062" points="652" swimtime="00:01:59.98" resultid="4085" heatid="4807" lane="2" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:04.10" />
                    <SPLIT distance="150" swimtime="00:01:32.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3945" number="1" />
                    <RELAYPOSITION athleteid="4024" number="2" />
                    <RELAYPOSITION athleteid="3926" number="3" />
                    <RELAYPOSITION athleteid="4064" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:50.00" eventid="2224" heatid="4810" lane="2" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5541" nation="GER" region="02" clubid="2503" name="SG Nordoberpfalz">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Kathrin" gender="F" lastname="Bachmeier" nation="GER" license="262269" athleteid="2504">
              <RESULTS>
                <RESULT eventid="1059" points="554" swimtime="00:01:01.98" resultid="2505" heatid="4669" lane="6" entrytime="00:01:02.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="425" swimtime="00:00:38.29" resultid="2506" heatid="4687" lane="5" entrytime="00:00:37.81" />
                <RESULT eventid="1785" points="406" swimtime="00:01:14.31" resultid="2507" heatid="4718" lane="5" entrytime="00:01:13.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="461" swimtime="00:01:13.35" resultid="2508" heatid="4730" lane="4" entrytime="00:01:13.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="528" swimtime="00:04:50.07" resultid="2509" heatid="4760" lane="2" entrytime="00:04:51.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:06.66" />
                    <SPLIT distance="150" swimtime="00:01:42.93" />
                    <SPLIT distance="200" swimtime="00:02:19.65" />
                    <SPLIT distance="250" swimtime="00:02:56.52" />
                    <SPLIT distance="300" swimtime="00:03:34.75" />
                    <SPLIT distance="350" swimtime="00:04:12.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:19.46" eventid="1978" heatid="4831" lane="1" />
                <ENTRY entrytime="00:02:39.19" eventid="2055" heatid="4897" lane="6" />
                <ENTRY entrytime="00:00:29.16" eventid="2082" heatid="4916" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lukas" gender="M" lastname="Bachmeier" nation="GER" license="210544" athleteid="2513">
              <RESULTS>
                <RESULT eventid="1763" points="417" swimtime="00:01:14.43" resultid="2514" heatid="4698" lane="1" entrytime="00:01:11.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="408" swimtime="00:02:27.73" resultid="2515" heatid="4751" lane="4" entrytime="00:02:21.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:11.12" />
                    <SPLIT distance="150" swimtime="00:01:52.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.73" eventid="1985" heatid="4843" lane="6" />
                <ENTRY entrytime="00:02:36.66" eventid="2089" heatid="4926" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Viktoria" gender="F" lastname="Bogner" nation="GER" license="287903" athleteid="2518">
              <RESULTS>
                <RESULT eventid="1059" points="485" swimtime="00:01:04.77" resultid="2519" heatid="4666" lane="6" entrytime="00:01:03.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="408" swimtime="00:00:38.82" resultid="2520" heatid="4687" lane="3" entrytime="00:00:37.54" />
                <RESULT eventid="1799" points="422" swimtime="00:01:15.53" resultid="2521" heatid="4729" lane="6" entrytime="00:01:14.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:20.52" eventid="1978" heatid="4830" lane="1" />
                <ENTRY entrytime="00:01:20.41" eventid="1992" heatid="4851" lane="4" />
                <ENTRY entrytime="00:00:29.74" eventid="2082" heatid="4914" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4305" nation="GER" region="02" clubid="3458" name="SG Oberland T.-I.-P. Penzberg">
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Florian" gender="M" lastname="De Witte" nation="GER" license="307167" athleteid="3459">
              <RESULTS>
                <RESULT eventid="1749" points="490" swimtime="00:02:06.03" resultid="3460" heatid="4679" lane="3" entrytime="00:02:04.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="100" swimtime="00:01:01.44" />
                    <SPLIT distance="150" swimtime="00:01:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="514" swimtime="00:01:00.46" resultid="3461" heatid="4712" lane="2" entrytime="00:01:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:15.83" eventid="2041" heatid="4894" lane="1" />
                <ENTRY entrytime="00:00:27.53" eventid="2103" heatid="4943" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Manuel" gender="M" lastname="Genster" nation="GER" license="240652" athleteid="3464">
              <RESULTS>
                <RESULT eventid="1749" points="636" swimtime="00:01:55.50" resultid="3465" heatid="4684" lane="5" entrytime="00:01:55.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                    <SPLIT distance="100" swimtime="00:00:55.58" />
                    <SPLIT distance="150" swimtime="00:01:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="623" swimtime="00:00:56.69" resultid="3466" heatid="4716" lane="3" entrytime="00:00:55.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="566" swimtime="00:00:24.48" resultid="3467" heatid="4775" lane="5" entrytime="00:00:24.05" />
                <RESULT eventid="1898" points="660" swimtime="00:00:55.63" resultid="5454" heatid="4717" lane="4" entrytime="00:00:56.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.15" eventid="1971" heatid="4826" lane="5" />
                <ENTRY entrytime="00:00:25.41" eventid="2103" heatid="4946" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Jakob" gender="M" lastname="Hoehler" nation="GER" license="246021" athleteid="3470">
              <RESULTS>
                <RESULT eventid="1763" points="470" swimtime="00:01:11.48" resultid="3471" heatid="4698" lane="3" entrytime="00:01:10.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.24" eventid="1985" heatid="4843" lane="3" />
                <ENTRY entrytime="00:02:35.80" eventid="2089" heatid="4927" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Philipp" gender="M" lastname="Kirchner" nation="GER" license="131299" athleteid="3474">
              <RESULTS>
                <RESULT eventid="1806" points="516" swimtime="00:00:27.69" resultid="3475" heatid="4743" lane="2" entrytime="00:00:27.87" />
                <RESULT eventid="1848" points="529" swimtime="00:02:10.54" resultid="3476" heatid="4789" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="150" swimtime="00:01:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1912" points="524" swimtime="00:00:27.56" resultid="5411" heatid="5417" lane="3" entrytime="00:00:27.69" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.65" eventid="2013" heatid="4871" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Martina Edda" gender="F" lastname="Lickel" nation="GER" license="284991" athleteid="3478">
              <RESULTS>
                <RESULT eventid="1059" points="594" swimtime="00:01:00.56" resultid="3479" heatid="4671" lane="3" entrytime="00:01:00.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="536" swimtime="00:01:07.73" resultid="3480" heatid="4723" lane="6" entrytime="00:01:08.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="606" swimtime="00:01:00.13" resultid="5329" heatid="5317" lane="6" entrytime="00:01:00.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:14.37" eventid="1978" heatid="4834" lane="5" />
                <ENTRY entrytime="00:00:32.21" eventid="2034" heatid="4887" lane="6" />
                <ENTRY entrytime="00:00:27.82" eventid="2082" heatid="4923" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Jonathan" gender="M" lastname="Schottenheim" nation="GER" license="306550" athleteid="3484">
              <RESULTS>
                <RESULT eventid="1763" points="439" swimtime="00:01:13.15" resultid="3485" heatid="4697" lane="2" entrytime="00:01:12.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.33" eventid="1985" heatid="4843" lane="4" />
                <ENTRY entrytime="00:02:38.72" eventid="2089" heatid="4926" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Sebastian" gender="M" lastname="Sonnenstuhl" nation="GER" license="226790" athleteid="3488">
              <RESULTS>
                <RESULT eventid="1820" points="458" swimtime="00:02:22.17" resultid="3489" heatid="4752" lane="3" entrytime="00:02:17.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:07.11" />
                    <SPLIT distance="150" swimtime="00:01:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="483" swimtime="00:00:25.82" resultid="3490" heatid="4773" lane="5" entrytime="00:00:25.03" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.22" eventid="1971" heatid="4820" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="543" swimtime="00:01:50.90" resultid="3492" heatid="4806" lane="6" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                    <SPLIT distance="100" swimtime="00:00:59.99" />
                    <SPLIT distance="150" swimtime="00:01:25.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3474" number="1" />
                    <RELAYPOSITION athleteid="3470" number="2" reactiontime="+46" />
                    <RELAYPOSITION athleteid="3464" number="3" reactiontime="+48" />
                    <RELAYPOSITION athleteid="3488" number="4" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6621" nation="GER" region="02" clubid="4242" name="SG Rödental">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Selina" gender="F" lastname="Jenke" nation="GER" license="265832" athleteid="4250">
              <RESULTS>
                <RESULT eventid="1059" points="556" swimtime="00:01:01.89" resultid="4251" heatid="4672" lane="6" entrytime="00:01:00.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="495" swimtime="00:00:30.80" resultid="4252" heatid="4798" lane="2" entrytime="00:00:30.77" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.88" eventid="2034" heatid="4886" lane="1" />
                <ENTRY entrytime="00:00:27.70" eventid="2082" heatid="4921" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Danielle" gender="F" lastname="Schuller" nation="GER" license="183972" athleteid="4255">
              <RESULTS>
                <RESULT eventid="1756" points="579" swimtime="00:00:34.54" resultid="4256" heatid="4691" lane="3" entrytime="00:00:35.43" />
                <RESULT eventid="1799" points="530" swimtime="00:01:10.02" resultid="4257" heatid="4735" lane="1" entrytime="00:01:11.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1877" points="594" swimtime="00:00:34.25" resultid="5353" heatid="5355" lane="1" entrytime="00:00:34.54" />
                <RESULT eventid="1919" points="529" swimtime="00:01:10.04" resultid="5400" heatid="5404" lane="2" entrytime="00:01:10.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:15.48" eventid="1992" heatid="4856" lane="2" />
                <ENTRY entrytime="00:00:28.59" eventid="2082" heatid="4918" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Maike" gender="F" lastname="Schuller" nation="GER" license="183954" athleteid="4260">
              <RESULTS>
                <RESULT eventid="1059" points="489" swimtime="00:01:04.61" resultid="4261" heatid="4663" lane="3" entrytime="00:01:04.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="496" swimtime="00:04:56.24" resultid="4262" heatid="4760" lane="1" entrytime="00:04:52.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                    <SPLIT distance="150" swimtime="00:01:45.16" />
                    <SPLIT distance="200" swimtime="00:02:23.40" />
                    <SPLIT distance="250" swimtime="00:03:01.72" />
                    <SPLIT distance="300" swimtime="00:03:40.14" />
                    <SPLIT distance="350" swimtime="00:04:19.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:20.57" eventid="1978" heatid="4830" lane="6" />
                <ENTRY entrytime="00:02:38.11" eventid="2055" heatid="4898" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.00" eventid="2224" heatid="4810" lane="6" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6423" nation="GER" region="02" clubid="2906" name="SG Stadtwerke München">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Sara" gender="F" lastname="Aringsmann" nation="GER" license="305291" athleteid="2922">
              <RESULTS>
                <RESULT eventid="1059" points="579" swimtime="00:01:01.08" resultid="2923" heatid="4667" lane="4" entrytime="00:01:02.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="602" swimtime="00:00:34.09" resultid="2924" heatid="4693" lane="1" entrytime="00:00:34.69" />
                <RESULT eventid="1841" points="602" swimtime="00:02:39.32" resultid="2925" heatid="4782" lane="5" entrytime="00:02:45.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:01:17.13" />
                    <SPLIT distance="150" swimtime="00:01:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1877" points="579" swimtime="00:00:34.55" resultid="5349" heatid="5355" lane="3" entrytime="00:00:34.09" />
                <RESULT eventid="1954" points="604" swimtime="00:02:39.15" resultid="5482" heatid="4785" lane="5" entrytime="00:02:39.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="150" swimtime="00:01:57.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:16.31" eventid="1992" heatid="4855" lane="1" />
                <ENTRY entrytime="00:02:31.62" eventid="2055" heatid="4903" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Yael" gender="M" lastname="Balz" nation="GER" license="318639" athleteid="2928">
              <RESULTS>
                <RESULT eventid="1792" points="608" swimtime="00:16:40.65" resultid="2929" heatid="4726" lane="3" entrytime="00:17:11.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="100" swimtime="00:01:01.66" />
                    <SPLIT distance="150" swimtime="00:01:35.33" />
                    <SPLIT distance="200" swimtime="00:02:08.84" />
                    <SPLIT distance="250" swimtime="00:02:42.47" />
                    <SPLIT distance="300" swimtime="00:03:16.39" />
                    <SPLIT distance="350" swimtime="00:03:50.38" />
                    <SPLIT distance="400" swimtime="00:04:24.08" />
                    <SPLIT distance="450" swimtime="00:04:58.19" />
                    <SPLIT distance="500" swimtime="00:05:32.19" />
                    <SPLIT distance="550" swimtime="00:06:05.51" />
                    <SPLIT distance="600" swimtime="00:06:39.44" />
                    <SPLIT distance="650" swimtime="00:07:13.20" />
                    <SPLIT distance="700" swimtime="00:07:47.03" />
                    <SPLIT distance="750" swimtime="00:08:21.12" />
                    <SPLIT distance="800" swimtime="00:08:54.94" />
                    <SPLIT distance="850" swimtime="00:09:28.76" />
                    <SPLIT distance="900" swimtime="00:10:01.92" />
                    <SPLIT distance="950" swimtime="00:10:35.23" />
                    <SPLIT distance="1000" swimtime="00:11:08.52" />
                    <SPLIT distance="1050" swimtime="00:11:42.08" />
                    <SPLIT distance="1100" swimtime="00:12:16.38" />
                    <SPLIT distance="1150" swimtime="00:12:49.75" />
                    <SPLIT distance="1200" swimtime="00:13:23.33" />
                    <SPLIT distance="1250" swimtime="00:13:56.70" />
                    <SPLIT distance="1300" swimtime="00:14:30.07" />
                    <SPLIT distance="1350" swimtime="00:15:03.57" />
                    <SPLIT distance="1400" swimtime="00:15:36.66" />
                    <SPLIT distance="1450" swimtime="00:16:09.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="418" swimtime="00:02:26.58" resultid="2930" heatid="4749" lane="2" entrytime="00:02:28.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="100" swimtime="00:01:11.11" />
                    <SPLIT distance="150" swimtime="00:01:54.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:15.37" eventid="2075" heatid="4910" lane="5" />
                <ENTRY entrytime="00:08:45.30" eventid="2168" heatid="4808" lane="5">
                  <MEETINFO qualificationtime="00:08:45.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Johanna" gender="F" lastname="Bander" nation="GER" license="281505" athleteid="2933">
              <RESULTS>
                <RESULT eventid="1827" points="540" swimtime="00:04:47.94" resultid="2934" heatid="4760" lane="3" entrytime="00:04:49.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:06.35" />
                    <SPLIT distance="150" swimtime="00:01:42.93" />
                    <SPLIT distance="200" swimtime="00:02:19.85" />
                    <SPLIT distance="250" swimtime="00:02:56.83" />
                    <SPLIT distance="300" swimtime="00:03:34.11" />
                    <SPLIT distance="350" swimtime="00:04:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="445" swimtime="00:00:31.91" resultid="2935" heatid="4795" lane="5" entrytime="00:00:31.74" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:22.21" eventid="1992" heatid="4850" lane="3" />
                <ENTRY entrytime="00:02:35.43" eventid="2055" heatid="4899" lane="3" />
                <ENTRY entrytime="00:00:29.07" eventid="2082" heatid="4916" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Janina" gender="F" lastname="Banse" nation="GER" license="234213" athleteid="2939">
              <RESULTS>
                <RESULT eventid="1059" points="637" swimtime="00:00:59.15" resultid="2940" heatid="4674" lane="4" entrytime="00:00:58.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1813" points="557" swimtime="00:02:25.36" resultid="2941" heatid="4747" lane="3" entrytime="00:02:17.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:10.06" />
                    <SPLIT distance="150" swimtime="00:01:48.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="690" swimtime="00:04:25.37" resultid="2942" heatid="4764" lane="4" entrytime="00:04:22.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:05.26" />
                    <SPLIT distance="150" swimtime="00:01:39.45" />
                    <SPLIT distance="200" swimtime="00:02:13.87" />
                    <SPLIT distance="250" swimtime="00:02:47.71" />
                    <SPLIT distance="300" swimtime="00:03:21.29" />
                    <SPLIT distance="350" swimtime="00:03:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="640" swimtime="00:00:59.05" resultid="5320" heatid="4675" lane="2" entrytime="00:00:59.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1933" points="569" swimtime="00:02:24.34" resultid="5422" heatid="4748" lane="1" entrytime="00:02:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:48.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:06.12" eventid="1978" heatid="4838" lane="4" />
                <ENTRY entrytime="00:01:04.11" eventid="2006" heatid="4866" lane="4" />
                <ENTRY entrytime="00:00:27.11" eventid="2082" heatid="4921" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Pascal" gender="M" lastname="Borchardt" nation="GER" license="287497" athleteid="2951">
              <RESULTS>
                <RESULT eventid="1749" points="466" swimtime="00:02:08.15" resultid="2952" heatid="4680" lane="4" entrytime="00:02:02.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="100" swimtime="00:01:00.85" />
                    <SPLIT distance="150" swimtime="00:01:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="492" swimtime="00:01:01.32" resultid="2953" heatid="4711" lane="4" entrytime="00:01:02.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="500" swimtime="00:00:25.52" resultid="2954" heatid="4772" lane="1" entrytime="00:00:25.42" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.51" eventid="1971" heatid="4821" lane="4" />
                <ENTRY entrytime="00:00:34.00" eventid="1985" heatid="4841" lane="3" />
                <ENTRY entrytime="00:01:08.46" eventid="2027" heatid="4877" lane="4" />
                <ENTRY entrytime="00:00:27.68" eventid="2103" heatid="4943" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Paulina" gender="F" lastname="Böger" nation="GER" license="202939" athleteid="2946">
              <RESULTS>
                <RESULT eventid="1756" points="633" swimtime="00:00:33.54" resultid="2947" heatid="4692" lane="4" entrytime="00:00:33.55" />
                <RESULT eventid="1841" points="598" swimtime="00:02:39.66" resultid="2948" heatid="4782" lane="4" entrytime="00:02:40.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:17.59" />
                    <SPLIT distance="150" swimtime="00:01:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1877" points="639" swimtime="00:00:33.42" resultid="5345" heatid="4695" lane="2" entrytime="00:00:33.54" />
                <RESULT eventid="1954" points="568" swimtime="00:02:42.45" resultid="5483" heatid="4785" lane="1" entrytime="00:02:39.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:18.73" />
                    <SPLIT distance="150" swimtime="00:02:00.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:13.38" eventid="1992" heatid="4856" lane="4" />
                <ENTRY entrytime="00:02:14.15" eventid="2096" heatid="4937" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lisa Marie" gender="F" lastname="Börnigen" nation="GER" license="267312" athleteid="2959">
              <RESULTS>
                <RESULT eventid="1059" points="611" swimtime="00:00:59.99" resultid="2960" heatid="4673" lane="6" entrytime="00:01:00.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1771" points="571" swimtime="00:05:12.62" resultid="2961" heatid="4708" lane="6" entrytime="00:05:14.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:49.80" />
                    <SPLIT distance="200" swimtime="00:02:29.60" />
                    <SPLIT distance="250" swimtime="00:03:15.38" />
                    <SPLIT distance="300" swimtime="00:04:01.88" />
                    <SPLIT distance="350" swimtime="00:04:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1813" points="505" swimtime="00:02:30.16" resultid="2962" heatid="4745" lane="5" entrytime="00:02:31.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:50.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="614" swimtime="00:00:59.87" resultid="5327" heatid="5317" lane="5" entrytime="00:00:59.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1933" points="536" swimtime="00:02:27.23" resultid="5426" heatid="5429" lane="2" entrytime="00:02:30.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:08.62" />
                    <SPLIT distance="150" swimtime="00:01:47.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:10:07.84" eventid="2020" status="RJC">
                  <MEETINFO qualificationtime="00:10:07.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.13" eventid="2096" heatid="4934" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Benjamin" gender="M" lastname="Campbell-James" nation="GER" license="376054" athleteid="2965">
              <RESULTS>
                <RESULT eventid="1778" points="474" swimtime="00:01:02.12" resultid="2966" heatid="4710" lane="1" entrytime="00:01:03.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="534" swimtime="00:02:15.11" resultid="2967" heatid="4753" lane="4" entrytime="00:02:14.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                    <SPLIT distance="100" swimtime="00:01:02.71" />
                    <SPLIT distance="150" swimtime="00:01:44.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="565" swimtime="00:02:07.71" resultid="2968" heatid="4790" lane="3" entrytime="00:02:07.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="100" swimtime="00:01:02.90" />
                    <SPLIT distance="150" swimtime="00:01:35.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="577" swimtime="00:02:06.83" resultid="5492" heatid="4792" lane="3" entrytime="00:02:07.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.00" />
                    <SPLIT distance="100" swimtime="00:01:02.45" />
                    <SPLIT distance="150" swimtime="00:01:35.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.12" eventid="1971" heatid="4822" lane="3" />
                <ENTRY entrytime="00:01:00.98" eventid="2013" heatid="4873" lane="5" />
                <ENTRY entrytime="00:04:18.09" eventid="2075" heatid="4910" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Elena" gender="F" lastname="Czeschner" nation="GER" license="183021" athleteid="2972">
              <RESULTS>
                <RESULT eventid="1059" points="617" swimtime="00:00:59.79" resultid="2973" heatid="4672" lane="3" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="578" swimtime="00:00:29.26" resultid="2974" heatid="4801" lane="3" entrytime="00:00:27.90" />
                <RESULT eventid="1940" points="585" swimtime="00:00:29.15" resultid="5509" heatid="4802" lane="1" entrytime="00:00:29.26" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:02.00" eventid="2006" heatid="4867" lane="3" />
                <ENTRY entrytime="00:00:26.31" eventid="2082" heatid="4923" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Henning" gender="M" lastname="Dörries" nation="GER" license="220261" athleteid="2977">
              <RESULTS>
                <RESULT eventid="1749" points="605" swimtime="00:01:57.45" resultid="2978" heatid="4685" lane="5" entrytime="00:01:55.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                    <SPLIT distance="100" swimtime="00:00:56.90" />
                    <SPLIT distance="150" swimtime="00:01:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1792" points="683" swimtime="00:16:02.75" resultid="2979" heatid="4727" lane="4" entrytime="00:16:06.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:32.30" />
                    <SPLIT distance="200" swimtime="00:02:04.38" />
                    <SPLIT distance="250" swimtime="00:02:36.36" />
                    <SPLIT distance="300" swimtime="00:03:08.36" />
                    <SPLIT distance="350" swimtime="00:03:40.28" />
                    <SPLIT distance="400" swimtime="00:04:12.48" />
                    <SPLIT distance="450" swimtime="00:04:45.07" />
                    <SPLIT distance="500" swimtime="00:05:17.61" />
                    <SPLIT distance="550" swimtime="00:05:50.08" />
                    <SPLIT distance="600" swimtime="00:06:22.30" />
                    <SPLIT distance="650" swimtime="00:06:54.84" />
                    <SPLIT distance="700" swimtime="00:07:26.84" />
                    <SPLIT distance="750" swimtime="00:07:59.51" />
                    <SPLIT distance="800" swimtime="00:08:31.92" />
                    <SPLIT distance="850" swimtime="00:09:04.86" />
                    <SPLIT distance="900" swimtime="00:09:37.31" />
                    <SPLIT distance="950" swimtime="00:10:09.85" />
                    <SPLIT distance="1000" swimtime="00:10:42.18" />
                    <SPLIT distance="1050" swimtime="00:11:14.70" />
                    <SPLIT distance="1100" swimtime="00:11:47.04" />
                    <SPLIT distance="1150" swimtime="00:12:19.41" />
                    <SPLIT distance="1200" swimtime="00:12:51.77" />
                    <SPLIT distance="1250" swimtime="00:13:24.19" />
                    <SPLIT distance="1300" swimtime="00:13:56.18" />
                    <SPLIT distance="1350" swimtime="00:14:28.21" />
                    <SPLIT distance="1400" swimtime="00:15:00.54" />
                    <SPLIT distance="1450" swimtime="00:15:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="507" swimtime="00:00:25.40" resultid="2980" heatid="4772" lane="2" entrytime="00:00:25.32" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:40.51" eventid="1999" heatid="4862" lane="6" />
                <ENTRY entrytime="00:01:03.55" eventid="2027" heatid="4878" lane="3" />
                <ENTRY entrytime="00:04:06.47" eventid="2075" heatid="4911" lane="3" />
                <ENTRY entrytime="00:08:29.14" eventid="2168" heatid="4809" lane="2">
                  <MEETINFO qualificationtime="00:08:29.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Anastasia" gender="F" lastname="Eftimova" nation="GER" license="323701" athleteid="2985">
              <RESULTS>
                <RESULT eventid="1059" points="476" swimtime="00:01:05.19" resultid="2986" heatid="4662" lane="5" entrytime="00:01:05.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="465" swimtime="00:00:37.16" resultid="2987" heatid="4689" lane="1" entrytime="00:00:37.02" />
                <RESULT eventid="1841" points="433" swimtime="00:02:57.81" resultid="2988" heatid="4779" lane="2" entrytime="00:02:57.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:25.30" />
                    <SPLIT distance="150" swimtime="00:02:11.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:20.04" eventid="1992" heatid="4852" lane="6" />
                <ENTRY entrytime="00:00:29.74" eventid="2082" heatid="4914" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Veronika" gender="F" lastname="Ehrenbauer" nation="GER" license="106748" athleteid="2991">
              <RESULTS>
                <RESULT eventid="1785" points="593" swimtime="00:01:05.48" resultid="2992" heatid="4724" lane="3" entrytime="00:01:01.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="598" swimtime="00:01:07.24" resultid="2993" heatid="4736" lane="3" entrytime="00:01:02.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="654" swimtime="00:00:28.08" resultid="2994" heatid="4961" lane="3" entrytime="00:00:27.18" />
                <RESULT eventid="1891" points="665" swimtime="00:01:03.02" resultid="5382" heatid="4725" lane="5" entrytime="00:01:05.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1919" points="663" swimtime="00:01:04.99" resultid="5395" heatid="4737" lane="5" entrytime="00:01:07.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="662" swimtime="00:00:27.96" resultid="5505" heatid="4802" lane="3" entrytime="00:00:28.08" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Konrad" gender="M" lastname="Fleckenstein" nation="GER" license="247730" athleteid="2995">
              <RESULTS>
                <RESULT eventid="1749" points="511" swimtime="00:02:04.22" resultid="2996" heatid="4681" lane="5" entrytime="00:02:02.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                    <SPLIT distance="100" swimtime="00:01:00.06" />
                    <SPLIT distance="150" swimtime="00:01:32.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="555" swimtime="00:00:58.92" resultid="2997" heatid="4715" lane="4" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="548" swimtime="00:00:24.75" resultid="2998" heatid="4776" lane="1" entrytime="00:00:24.44" />
                <RESULT eventid="1898" points="585" swimtime="00:00:57.90" resultid="5461" heatid="5465" lane="2" entrytime="00:00:58.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.33" eventid="1971" heatid="4823" lane="4" />
                <ENTRY entrytime="00:02:10.00" eventid="2041" heatid="4894" lane="2" />
                <ENTRY entrytime="00:00:25.50" eventid="2103" heatid="4946" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Rabea" gender="F" lastname="Gärtner" nation="GER" license="316345" athleteid="3002">
              <RESULTS>
                <RESULT eventid="1059" points="464" swimtime="00:01:05.74" resultid="3003" heatid="4662" lane="3" entrytime="00:01:04.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="444" swimtime="00:00:37.74" resultid="3004" heatid="4688" lane="5" entrytime="00:00:37.39" />
                <RESULT eventid="1799" points="440" swimtime="00:01:14.46" resultid="3005" heatid="4729" lane="3" entrytime="00:01:14.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="492" swimtime="00:02:50.43" resultid="3006" heatid="4781" lane="6" entrytime="00:02:51.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:01:22.21" />
                    <SPLIT distance="150" swimtime="00:02:06.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:20.08" eventid="1992" heatid="4851" lane="3" />
                <ENTRY entrytime="00:02:40.18" eventid="2055" heatid="4896" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Benno" gender="M" lastname="Hawe" nation="GER" license="68494" athleteid="3009">
              <RESULTS>
                <RESULT eventid="1763" points="647" swimtime="00:01:04.27" resultid="3010" heatid="4702" lane="4" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1884" points="642" swimtime="00:01:04.45" resultid="5362" heatid="5368" lane="3" entrytime="00:01:04.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.54" eventid="1985" heatid="4847" lane="2" />
                <ENTRY entrytime="00:02:15.00" eventid="2089" heatid="4929" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Anna" gender="F" lastname="Herbst" nation="GER" license="250303" athleteid="3013">
              <RESULTS>
                <RESULT eventid="1785" points="574" swimtime="00:01:06.21" resultid="3014" heatid="4723" lane="5" entrytime="00:01:05.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1813" points="500" swimtime="00:02:30.65" resultid="3015" heatid="4745" lane="2" entrytime="00:02:28.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:52.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="531" swimtime="00:00:30.09" resultid="3016" heatid="4961" lane="5" entrytime="00:00:29.53" />
                <RESULT eventid="1891" points="570" swimtime="00:01:06.35" resultid="5386" heatid="5391" lane="4" entrytime="00:01:06.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="556" swimtime="00:00:29.64" resultid="5514" heatid="5517" lane="5" entrytime="00:00:30.09" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="2006" heatid="4867" lane="2" />
                <ENTRY entrytime="00:00:31.72" eventid="2034" heatid="4889" lane="1" />
                <ENTRY entrytime="00:02:28.00" eventid="2055" heatid="4904" lane="1" />
                <ENTRY entrytime="00:02:27.29" eventid="2096" heatid="4936" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Anastasia" gender="F" lastname="Ismyrli" nation="GER" license="332675" athleteid="3021">
              <RESULTS>
                <RESULT eventid="1756" points="645" swimtime="00:00:33.33" resultid="3022" heatid="4693" lane="3" entrytime="00:00:32.71" />
                <RESULT eventid="1841" points="627" swimtime="00:02:37.17" resultid="3023" heatid="4784" lane="4" entrytime="00:02:38.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:01:56.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="512" swimtime="00:00:30.46" resultid="3024" heatid="4961" lane="6" entrytime="00:00:29.89" />
                <RESULT eventid="1877" points="635" swimtime="00:00:33.49" resultid="5344" heatid="4695" lane="4" entrytime="00:00:33.33" />
                <RESULT eventid="1954" points="607" swimtime="00:02:38.87" resultid="5480" heatid="4785" lane="4" entrytime="00:02:37.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:01:15.88" />
                    <SPLIT distance="150" swimtime="00:01:57.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:11.63" eventid="1992" heatid="4856" lane="3" />
                <ENTRY entrytime="00:01:05.72" eventid="2006" heatid="4865" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Sebastian" gender="M" lastname="Koller" nation="GER" license="184756" athleteid="3027">
              <RESULTS>
                <RESULT eventid="1763" points="620" swimtime="00:01:05.19" resultid="3028" heatid="4703" lane="2" entrytime="00:01:04.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="(Zeit: 17:26), Schwimmer hat bei der 50m Wende nicht mit beiden Händen gelichzeitig angeschlagen." eventid="1884" status="DSQ" swimtime="00:01:04.83" resultid="5367" heatid="5368" lane="6" entrytime="00:01:05.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.42" eventid="1985" heatid="4848" lane="2" />
                <ENTRY entrytime="00:02:16.45" eventid="2089" heatid="4928" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Stella" gender="F" lastname="Koltermann" nation="GER" license="245421" athleteid="3031">
              <RESULTS>
                <RESULT eventid="1785" status="DNS" swimtime="00:00:00.00" resultid="3032" heatid="4720" lane="3" entrytime="00:01:10.87" />
                <RESULT eventid="1855" status="DNS" swimtime="00:00:00.00" resultid="3033" heatid="4797" lane="6" entrytime="00:00:31.17" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:14.22" eventid="1978" heatid="4834" lane="2" />
                <ENTRY entrytime="00:00:28.28" eventid="2082" heatid="4920" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Victoria" gender="F" lastname="Kothny" nation="GER" license="274693" athleteid="3201">
              <RESULTS>
                <RESULT eventid="1059" points="546" swimtime="00:01:02.26" resultid="3202" heatid="4672" lane="1" entrytime="00:01:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="571" swimtime="00:01:06.31" resultid="3203" heatid="4722" lane="2" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="604" swimtime="00:04:37.40" resultid="3204" heatid="4762" lane="1" entrytime="00:04:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:06.03" />
                    <SPLIT distance="150" swimtime="00:01:41.34" />
                    <SPLIT distance="200" swimtime="00:02:17.36" />
                    <SPLIT distance="250" swimtime="00:02:52.65" />
                    <SPLIT distance="300" swimtime="00:03:28.07" />
                    <SPLIT distance="350" swimtime="00:04:03.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1891" points="587" swimtime="00:01:05.69" resultid="5387" heatid="5391" lane="2" entrytime="00:01:06.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:12.50" eventid="1978" heatid="4835" lane="2" />
                <ENTRY entrytime="00:00:30.41" eventid="2034" heatid="4889" lane="4" />
                <ENTRY entrytime="00:02:21.88" eventid="2096" heatid="4937" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Robert" gender="M" lastname="Könneker" nation="GER" license="75201" athleteid="3036">
              <RESULTS>
                <RESULT eventid="1806" points="705" swimtime="00:00:24.96" resultid="3037" heatid="4743" lane="3" entrytime="00:00:24.49" />
                <RESULT eventid="1834" points="748" swimtime="00:00:22.31" resultid="3038" heatid="4776" lane="3" entrytime="00:00:22.91" />
                <RESULT eventid="1912" points="714" swimtime="00:00:24.85" resultid="5405" heatid="4744" lane="3" entrytime="00:00:24.96" />
                <RESULT eventid="1947" points="744" swimtime="00:00:22.35" resultid="5466" heatid="4778" lane="3" entrytime="00:00:22.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Amelie" gender="F" lastname="Liesenfeld" nation="GER" license="301144" athleteid="3039">
              <RESULTS>
                <RESULT eventid="1756" points="530" swimtime="00:00:35.57" resultid="3040" heatid="4690" lane="5" entrytime="00:00:36.23" />
                <RESULT eventid="1771" points="472" swimtime="00:05:33.18" resultid="3041" heatid="4705" lane="3" entrytime="00:05:39.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="150" swimtime="00:02:04.49" />
                    <SPLIT distance="200" swimtime="00:02:45.89" />
                    <SPLIT distance="250" swimtime="00:03:30.79" />
                    <SPLIT distance="300" swimtime="00:04:16.18" />
                    <SPLIT distance="350" swimtime="00:04:55.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="468" swimtime="00:01:12.94" resultid="3042" heatid="4729" lane="4" entrytime="00:01:14.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="529" swimtime="00:02:46.29" resultid="3043" heatid="4782" lane="1" entrytime="00:02:46.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:04.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:17.21" eventid="1992" heatid="4854" lane="2" />
                <ENTRY entrytime="00:02:38.64" eventid="2055" heatid="4897" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Luisa" gender="F" lastname="Liesenfeld" nation="GER" license="297730" athleteid="3046">
              <RESULTS>
                <RESULT eventid="1059" points="517" swimtime="00:01:03.40" resultid="3047" heatid="4663" lane="1" entrytime="00:01:04.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="553" swimtime="00:04:45.61" resultid="3048" heatid="4762" lane="6" entrytime="00:04:42.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                    <SPLIT distance="150" swimtime="00:01:43.68" />
                    <SPLIT distance="200" swimtime="00:02:20.30" />
                    <SPLIT distance="250" swimtime="00:02:57.12" />
                    <SPLIT distance="300" swimtime="00:03:33.90" />
                    <SPLIT distance="350" swimtime="00:04:10.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="561" swimtime="00:18:34.86" resultid="3049" heatid="4803" lane="4" entrytime="00:18:42.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                    <SPLIT distance="100" swimtime="00:01:08.24" />
                    <SPLIT distance="150" swimtime="00:01:44.73" />
                    <SPLIT distance="200" swimtime="00:02:21.65" />
                    <SPLIT distance="250" swimtime="00:02:58.85" />
                    <SPLIT distance="300" swimtime="00:03:35.82" />
                    <SPLIT distance="350" swimtime="00:04:13.09" />
                    <SPLIT distance="400" swimtime="00:04:50.28" />
                    <SPLIT distance="450" swimtime="00:05:27.65" />
                    <SPLIT distance="500" swimtime="00:06:05.31" />
                    <SPLIT distance="550" swimtime="00:06:42.57" />
                    <SPLIT distance="600" swimtime="00:07:19.94" />
                    <SPLIT distance="650" swimtime="00:07:57.58" />
                    <SPLIT distance="700" swimtime="00:08:35.50" />
                    <SPLIT distance="750" swimtime="00:09:13.11" />
                    <SPLIT distance="800" swimtime="00:09:50.98" />
                    <SPLIT distance="850" swimtime="00:10:28.57" />
                    <SPLIT distance="900" swimtime="00:11:06.54" />
                    <SPLIT distance="950" swimtime="00:11:44.15" />
                    <SPLIT distance="1000" swimtime="00:12:21.55" />
                    <SPLIT distance="1050" swimtime="00:12:59.67" />
                    <SPLIT distance="1100" swimtime="00:13:37.79" />
                    <SPLIT distance="1150" swimtime="00:14:15.10" />
                    <SPLIT distance="1200" swimtime="00:14:53.12" />
                    <SPLIT distance="1250" swimtime="00:15:30.76" />
                    <SPLIT distance="1300" swimtime="00:16:08.55" />
                    <SPLIT distance="1350" swimtime="00:16:45.51" />
                    <SPLIT distance="1400" swimtime="00:17:22.48" />
                    <SPLIT distance="1450" swimtime="00:17:59.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:16.10" eventid="1978" heatid="4832" lane="3" />
                <ENTRY entrytime="00:09:48.60" eventid="2020" heatid="4875" lane="2">
                  <MEETINFO qualificationtime="00:09:48.60" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Anna" gender="F" lastname="Metzler" nation="GER" license="278615" athleteid="3058">
              <RESULTS>
                <RESULT eventid="1059" points="630" swimtime="00:00:59.37" resultid="3059" heatid="4674" lane="1" entrytime="00:01:00.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="578" swimtime="00:01:06.04" resultid="3060" heatid="4724" lane="5" entrytime="00:01:05.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="616" swimtime="00:02:38.10" resultid="3061" heatid="4782" lane="2" entrytime="00:02:44.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.57" />
                    <SPLIT distance="100" swimtime="00:01:17.75" />
                    <SPLIT distance="150" swimtime="00:01:58.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="627" swimtime="00:00:59.45" resultid="5321" heatid="4675" lane="5" entrytime="00:00:59.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1891" points="550" swimtime="00:01:07.13" resultid="5384" heatid="4725" lane="6" entrytime="00:01:06.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:06.56" eventid="1978" heatid="4837" lane="4" />
                <ENTRY entrytime="00:01:06.36" eventid="2006" heatid="4866" lane="5" />
                <ENTRY entrytime="00:02:22.81" eventid="2055" heatid="4902" lane="4" />
                <ENTRY entrytime="00:02:23.00" eventid="2096" heatid="4936" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Andreas" gender="M" lastname="März" nation="GER" license="301258" athleteid="3052">
              <RESULTS>
                <RESULT eventid="1792" points="602" swimtime="00:16:43.94" resultid="3053" heatid="4726" lane="2" entrytime="00:17:51.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:02.46" />
                    <SPLIT distance="150" swimtime="00:01:35.75" />
                    <SPLIT distance="200" swimtime="00:02:09.28" />
                    <SPLIT distance="250" swimtime="00:02:42.67" />
                    <SPLIT distance="300" swimtime="00:03:16.67" />
                    <SPLIT distance="350" swimtime="00:03:50.51" />
                    <SPLIT distance="400" swimtime="00:04:24.35" />
                    <SPLIT distance="450" swimtime="00:04:58.55" />
                    <SPLIT distance="500" swimtime="00:05:31.88" />
                    <SPLIT distance="550" swimtime="00:06:05.62" />
                    <SPLIT distance="600" swimtime="00:06:39.54" />
                    <SPLIT distance="650" swimtime="00:07:13.53" />
                    <SPLIT distance="700" swimtime="00:07:47.12" />
                    <SPLIT distance="750" swimtime="00:08:21.44" />
                    <SPLIT distance="800" swimtime="00:08:54.94" />
                    <SPLIT distance="850" swimtime="00:09:29.09" />
                    <SPLIT distance="900" swimtime="00:10:02.44" />
                    <SPLIT distance="950" swimtime="00:10:36.26" />
                    <SPLIT distance="1000" swimtime="00:11:09.71" />
                    <SPLIT distance="1050" swimtime="00:11:43.13" />
                    <SPLIT distance="1100" swimtime="00:12:16.93" />
                    <SPLIT distance="1150" swimtime="00:12:50.90" />
                    <SPLIT distance="1200" swimtime="00:13:24.43" />
                    <SPLIT distance="1250" swimtime="00:13:57.66" />
                    <SPLIT distance="1300" swimtime="00:14:31.40" />
                    <SPLIT distance="1350" swimtime="00:15:05.05" />
                    <SPLIT distance="1400" swimtime="00:15:38.45" />
                    <SPLIT distance="1450" swimtime="00:16:11.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="512" swimtime="00:02:11.97" resultid="3054" heatid="4790" lane="1" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                    <SPLIT distance="150" swimtime="00:01:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="495" swimtime="00:02:13.51" resultid="5496" heatid="4792" lane="1" entrytime="00:02:11.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:05.56" />
                    <SPLIT distance="150" swimtime="00:01:40.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:50.04" eventid="1999" heatid="4861" lane="1" />
                <ENTRY entrytime="00:01:00.90" eventid="2013" heatid="4871" lane="2" />
                <ENTRY entrytime="00:02:40.53" eventid="2089" heatid="4925" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Mara" gender="F" lastname="Münsch" nation="GER" license="280574" athleteid="3066">
              <RESULTS>
                <RESULT eventid="1771" points="484" swimtime="00:05:30.34" resultid="3067" heatid="4706" lane="2" entrytime="00:05:32.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:02:00.31" />
                    <SPLIT distance="200" swimtime="00:02:41.23" />
                    <SPLIT distance="250" swimtime="00:03:28.03" />
                    <SPLIT distance="300" swimtime="00:04:16.50" />
                    <SPLIT distance="350" swimtime="00:04:53.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="441" swimtime="00:01:14.40" resultid="3068" heatid="4728" lane="5" entrytime="00:01:15.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="518" swimtime="00:04:52.01" resultid="3069" heatid="4760" lane="4" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:45.01" />
                    <SPLIT distance="200" swimtime="00:02:22.19" />
                    <SPLIT distance="250" swimtime="00:02:59.96" />
                    <SPLIT distance="300" swimtime="00:03:37.84" />
                    <SPLIT distance="350" swimtime="00:04:15.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:19.98" eventid="1978" heatid="4830" lane="3" />
                <ENTRY entrytime="00:02:38.79" eventid="2055" heatid="4897" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Max" gender="M" lastname="Nowosad" nation="GER" license="170324" athleteid="3072">
              <RESULTS>
                <RESULT eventid="1749" points="709" swimtime="00:01:51.42" resultid="3073" heatid="4685" lane="3" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                    <SPLIT distance="100" swimtime="00:00:54.63" />
                    <SPLIT distance="150" swimtime="00:01:23.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="659" swimtime="00:02:05.94" resultid="3074" heatid="4756" lane="4" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="100" swimtime="00:00:59.92" />
                    <SPLIT distance="150" swimtime="00:01:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="697" swimtime="00:02:03.63" resultid="5430" heatid="4757" lane="3" entrytime="00:02:05.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                    <SPLIT distance="100" swimtime="00:00:59.75" />
                    <SPLIT distance="150" swimtime="00:01:36.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:51.76" eventid="1971" heatid="4825" lane="4" />
                <ENTRY entrytime="00:02:05.00" eventid="2041" heatid="4893" lane="3" />
                <ENTRY entrytime="00:03:49.00" eventid="2075" heatid="4912" lane="4" />
                <ENTRY entrytime="NT" eventid="2168" status="RJC" />
                <ENTRY entrytime="00:01:51.42" eventid="1870" heatid="4686" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Christopher" gender="M" lastname="Richter" nation="GER" license="278786" athleteid="3079">
              <RESULTS>
                <RESULT eventid="1749" points="630" swimtime="00:01:55.86" resultid="3080" heatid="4683" lane="2" entrytime="00:01:54.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.99" />
                    <SPLIT distance="100" swimtime="00:00:56.73" />
                    <SPLIT distance="150" swimtime="00:01:27.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="524" swimtime="00:01:00.06" resultid="3081" heatid="4712" lane="5" entrytime="00:01:01.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="520" swimtime="00:00:25.18" resultid="3082" heatid="4772" lane="3" entrytime="00:00:25.16" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.44" eventid="1971" heatid="4825" lane="1" />
                <ENTRY entrytime="00:04:13.87" eventid="2075" heatid="4910" lane="2" />
                <ENTRY entrytime="00:08:40.79" eventid="2168" heatid="4808" lane="2">
                  <MEETINFO qualificationtime="00:08:39.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.86" eventid="1870" heatid="5342" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Felix" gender="M" lastname="Richtsfeld" nation="GER" license="223387" athleteid="3086">
              <RESULTS>
                <RESULT eventid="1749" points="674" swimtime="00:01:53.33" resultid="3087" heatid="4685" lane="1" entrytime="00:01:56.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                    <SPLIT distance="100" swimtime="00:00:55.99" />
                    <SPLIT distance="150" swimtime="00:01:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="587" swimtime="00:02:10.90" resultid="3088" heatid="4756" lane="6" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="100" swimtime="00:01:02.59" />
                    <SPLIT distance="150" swimtime="00:01:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="596" swimtime="00:02:10.23" resultid="5439" heatid="5442" lane="5" entrytime="00:02:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="100" swimtime="00:01:02.19" />
                    <SPLIT distance="150" swimtime="00:01:41.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.54" eventid="1971" heatid="4827" lane="6" />
                <ENTRY entrytime="00:04:03.00" eventid="2075" heatid="4912" lane="1" />
                <ENTRY entrytime="00:08:35.70" eventid="2168" heatid="4808" lane="4">
                  <MEETINFO qualificationtime="00:08:35.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.33" eventid="1870" heatid="4686" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Derik" gender="M" lastname="Rodrigues" nation="GER" license="245161" athleteid="3092">
              <RESULTS>
                <RESULT eventid="1749" points="554" swimtime="00:02:00.99" resultid="3093" heatid="4679" lane="4" entrytime="00:02:04.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                    <SPLIT distance="100" swimtime="00:00:57.75" />
                    <SPLIT distance="150" swimtime="00:01:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="556" swimtime="00:00:58.88" resultid="3094" heatid="4715" lane="5" entrytime="00:00:59.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="512" swimtime="00:02:16.96" resultid="3095" heatid="4752" lane="5" entrytime="00:02:19.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                    <SPLIT distance="100" swimtime="00:01:04.53" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1898" points="551" swimtime="00:00:59.06" resultid="5459" heatid="5465" lane="3" entrytime="00:00:58.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.00" eventid="1971" heatid="4818" lane="1" />
                <ENTRY entrytime="00:01:01.93" eventid="2013" heatid="4873" lane="1" />
                <ENTRY entrytime="00:02:10.00" eventid="2041" heatid="4892" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Aleksandar" gender="M" lastname="Savic" nation="GER" license="292599" athleteid="3099">
              <RESULTS>
                <RESULT eventid="1749" points="519" swimtime="00:02:03.61" resultid="3100" heatid="4679" lane="1" entrytime="00:02:05.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="100" swimtime="00:00:58.85" />
                    <SPLIT distance="150" swimtime="00:01:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="421" swimtime="00:01:04.63" resultid="3101" heatid="4711" lane="1" entrytime="00:01:02.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="501" swimtime="00:00:25.50" resultid="3102" heatid="4770" lane="5" entrytime="00:00:25.98" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.97" eventid="1971" heatid="4818" lane="2" />
                <ENTRY entrytime="00:01:06.50" eventid="2013" heatid="4869" lane="6" />
                <ENTRY entrytime="00:04:24.68" eventid="2075" heatid="4909" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Dajana" gender="F" lastname="Schlegel" nation="GER" license="158544" athleteid="3106">
              <RESULTS>
                <RESULT eventid="1059" points="575" swimtime="00:01:01.21" resultid="3107" heatid="4670" lane="2" entrytime="00:01:01.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="644" swimtime="00:01:03.72" resultid="3108" heatid="4722" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="692" swimtime="00:04:25.13" resultid="3109" heatid="4764" lane="1" entrytime="00:04:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:04.32" />
                    <SPLIT distance="150" swimtime="00:01:38.45" />
                    <SPLIT distance="200" swimtime="00:02:12.28" />
                    <SPLIT distance="250" swimtime="00:02:45.92" />
                    <SPLIT distance="300" swimtime="00:03:19.51" />
                    <SPLIT distance="350" swimtime="00:03:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1891" points="644" swimtime="00:01:03.71" resultid="5379" heatid="4725" lane="3" entrytime="00:01:03.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:11.00" eventid="1978" heatid="4837" lane="6" />
                <ENTRY entrytime="00:00:31.40" eventid="2034" heatid="4888" lane="5" />
                <ENTRY entrytime="00:02:28.00" eventid="2055" heatid="4903" lane="1" />
                <ENTRY entrytime="00:02:18.00" eventid="2096" heatid="4936" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Lisa Ava" gender="F" lastname="Schlüter" nation="GER" license="310203" athleteid="3114">
              <RESULTS>
                <RESULT eventid="1059" points="505" swimtime="00:01:03.92" resultid="3115" heatid="4666" lane="2" entrytime="00:01:03.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="421" swimtime="00:01:13.39" resultid="3116" heatid="4718" lane="2" entrytime="00:01:13.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="557" swimtime="00:18:37.26" resultid="3117" heatid="4803" lane="6" entrytime="00:19:00.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:44.71" />
                    <SPLIT distance="200" swimtime="00:02:21.82" />
                    <SPLIT distance="250" swimtime="00:02:59.06" />
                    <SPLIT distance="300" swimtime="00:03:36.36" />
                    <SPLIT distance="350" swimtime="00:04:13.95" />
                    <SPLIT distance="400" swimtime="00:04:51.62" />
                    <SPLIT distance="450" swimtime="00:05:29.39" />
                    <SPLIT distance="500" swimtime="00:06:07.08" />
                    <SPLIT distance="550" swimtime="00:06:44.93" />
                    <SPLIT distance="600" swimtime="00:07:22.68" />
                    <SPLIT distance="650" swimtime="00:08:00.58" />
                    <SPLIT distance="700" swimtime="00:08:38.42" />
                    <SPLIT distance="750" swimtime="00:09:16.22" />
                    <SPLIT distance="800" swimtime="00:09:54.05" />
                    <SPLIT distance="850" swimtime="00:10:31.76" />
                    <SPLIT distance="900" swimtime="00:11:09.24" />
                    <SPLIT distance="950" swimtime="00:11:46.87" />
                    <SPLIT distance="1000" swimtime="00:12:24.51" />
                    <SPLIT distance="1050" swimtime="00:13:02.07" />
                    <SPLIT distance="1100" swimtime="00:13:39.73" />
                    <SPLIT distance="1150" swimtime="00:14:17.34" />
                    <SPLIT distance="1200" swimtime="00:14:54.96" />
                    <SPLIT distance="1250" swimtime="00:15:32.83" />
                    <SPLIT distance="1300" swimtime="00:16:10.44" />
                    <SPLIT distance="1350" swimtime="00:16:47.94" />
                    <SPLIT distance="1400" swimtime="00:17:25.33" />
                    <SPLIT distance="1450" swimtime="00:18:02.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:15.09" eventid="1978" heatid="4834" lane="6" />
                <ENTRY entrytime="00:10:03.80" eventid="2020" status="RJC">
                  <MEETINFO qualificationtime="00:09:59.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.37" eventid="2096" heatid="4933" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Marc" gender="M" lastname="Schmid" nation="GER" license="186315" athleteid="3127">
              <RESULTS>
                <RESULT eventid="1763" points="685" swimtime="00:01:03.08" resultid="3128" heatid="4701" lane="4" entrytime="00:01:04.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="642" swimtime="00:02:07.08" resultid="3129" heatid="4755" lane="3" entrytime="00:02:04.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                    <SPLIT distance="100" swimtime="00:01:00.69" />
                    <SPLIT distance="150" swimtime="00:01:37.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="523" swimtime="00:02:11.04" resultid="3130" heatid="4791" lane="4" entrytime="00:02:09.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:01:03.85" />
                    <SPLIT distance="150" swimtime="00:01:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1884" points="689" swimtime="00:01:02.96" resultid="5358" heatid="4704" lane="2" entrytime="00:01:03.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="677" swimtime="00:02:04.82" resultid="5432" heatid="4757" lane="2" entrytime="00:02:07.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                    <SPLIT distance="100" swimtime="00:01:00.18" />
                    <SPLIT distance="150" swimtime="00:01:35.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:23.02" eventid="1999" heatid="4862" lane="3" />
                <ENTRY entrytime="00:02:04.67" eventid="2041" heatid="4894" lane="3" />
                <ENTRY entrytime="00:02:17.62" eventid="2089" heatid="4930" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Christoph" gender="M" lastname="Thade" nation="GER" license="132608" athleteid="3134">
              <RESULTS>
                <RESULT eventid="1749" points="524" swimtime="00:02:03.22" resultid="3135" heatid="4681" lane="4" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:00:59.38" />
                    <SPLIT distance="150" swimtime="00:01:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="506" swimtime="00:00:27.88" resultid="3136" heatid="4742" lane="3" entrytime="00:00:25.95" />
                <RESULT eventid="1834" points="569" swimtime="00:00:24.44" resultid="3137" heatid="4775" lane="3" entrytime="00:00:23.08" />
                <RESULT eventid="1912" points="511" swimtime="00:00:27.78" resultid="5413" heatid="5417" lane="2" entrytime="00:00:27.88" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:52.00" eventid="1971" heatid="4826" lane="2" />
                <ENTRY entrytime="00:00:57.68" eventid="2013" heatid="4872" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Titze" nation="GER" license="272986" athleteid="3140">
              <RESULTS>
                <RESULT eventid="1756" points="692" swimtime="00:00:32.56" resultid="3141" heatid="4694" lane="3" entrytime="00:00:32.56" />
                <RESULT eventid="1785" points="521" swimtime="00:01:08.38" resultid="3142" heatid="4722" lane="3" entrytime="00:01:04.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="622" swimtime="00:01:06.38" resultid="3143" heatid="4735" lane="3" entrytime="00:01:04.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="515" swimtime="00:00:30.41" resultid="3144" heatid="4801" lane="1" entrytime="00:00:29.74" />
                <RESULT eventid="1877" points="666" swimtime="00:00:32.97" resultid="5343" heatid="4695" lane="3" entrytime="00:00:32.56" />
                <RESULT eventid="1919" points="639" swimtime="00:01:05.76" resultid="5393" heatid="4737" lane="4" entrytime="00:01:06.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:12.72" eventid="1992" heatid="4855" lane="3" />
                <ENTRY entrytime="00:00:30.24" eventid="2034" heatid="4887" lane="3" />
                <ENTRY entrytime="00:02:22.39" eventid="2055" heatid="4903" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Sarah" gender="F" lastname="Vidic" nation="GER" license="290443" athleteid="3148">
              <RESULTS>
                <RESULT eventid="1771" points="541" swimtime="00:05:18.29" resultid="3149" heatid="4707" lane="6" entrytime="00:05:28.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:14.55" />
                    <SPLIT distance="150" swimtime="00:01:52.12" />
                    <SPLIT distance="200" swimtime="00:02:30.25" />
                    <SPLIT distance="250" swimtime="00:03:17.06" />
                    <SPLIT distance="300" swimtime="00:04:04.04" />
                    <SPLIT distance="350" swimtime="00:04:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="527" swimtime="00:01:08.12" resultid="3150" heatid="4723" lane="1" entrytime="00:01:07.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.32" eventid="2034" heatid="4886" lane="3" />
                <ENTRY entrytime="00:02:32.79" eventid="2055" heatid="4901" lane="4" />
                <ENTRY entrytime="00:02:24.13" eventid="2096" heatid="4937" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Grant" gender="M" lastname="Wasserman" nation="GER" license="374576" athleteid="3154">
              <RESULTS>
                <RESULT eventid="1749" points="537" swimtime="00:02:02.21" resultid="3155" heatid="4681" lane="6" entrytime="00:02:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="100" swimtime="00:00:59.87" />
                    <SPLIT distance="150" swimtime="00:01:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="451" swimtime="00:01:03.12" resultid="3156" heatid="4709" lane="4" entrytime="00:01:04.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="433" swimtime="00:00:29.36" resultid="3157" heatid="4742" lane="1" entrytime="00:00:28.88" />
                <RESULT eventid="1834" status="DNS" swimtime="00:00:00.00" resultid="3158" heatid="4773" lane="4" entrytime="00:00:24.95" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.50" eventid="1971" heatid="4821" lane="3" />
                <ENTRY entrytime="00:01:02.28" eventid="2013" heatid="4873" lane="6" />
                <ENTRY entrytime="00:04:27.29" eventid="2075" heatid="4908" lane="3" />
                <ENTRY entrytime="00:00:28.11" eventid="2103" heatid="4941" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Sebastian" gender="M" lastname="Wenk" nation="GER" license="182900" athleteid="3163">
              <RESULTS>
                <RESULT eventid="1749" points="601" swimtime="00:01:57.74" resultid="3164" heatid="4682" lane="2" entrytime="00:02:00.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                    <SPLIT distance="100" swimtime="00:00:57.88" />
                    <SPLIT distance="150" swimtime="00:01:28.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="527" swimtime="00:00:59.96" resultid="3165" heatid="4713" lane="1" entrytime="00:01:01.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1792" points="635" swimtime="00:16:26.64" resultid="3166" heatid="4727" lane="5" entrytime="00:16:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="100" swimtime="00:01:01.65" />
                    <SPLIT distance="150" swimtime="00:01:34.45" />
                    <SPLIT distance="200" swimtime="00:02:07.21" />
                    <SPLIT distance="250" swimtime="00:02:40.11" />
                    <SPLIT distance="300" swimtime="00:03:13.17" />
                    <SPLIT distance="350" swimtime="00:03:46.12" />
                    <SPLIT distance="400" swimtime="00:04:18.84" />
                    <SPLIT distance="450" swimtime="00:04:51.80" />
                    <SPLIT distance="500" swimtime="00:05:25.28" />
                    <SPLIT distance="550" swimtime="00:05:58.28" />
                    <SPLIT distance="600" swimtime="00:06:31.37" />
                    <SPLIT distance="650" swimtime="00:07:04.37" />
                    <SPLIT distance="700" swimtime="00:07:37.72" />
                    <SPLIT distance="750" swimtime="00:08:10.90" />
                    <SPLIT distance="800" swimtime="00:08:43.42" />
                    <SPLIT distance="850" swimtime="00:09:16.92" />
                    <SPLIT distance="900" swimtime="00:09:50.24" />
                    <SPLIT distance="950" swimtime="00:10:24.07" />
                    <SPLIT distance="1000" swimtime="00:10:57.65" />
                    <SPLIT distance="1050" swimtime="00:11:30.87" />
                    <SPLIT distance="1100" swimtime="00:12:04.50" />
                    <SPLIT distance="1150" swimtime="00:12:37.45" />
                    <SPLIT distance="1200" swimtime="00:13:10.21" />
                    <SPLIT distance="1250" swimtime="00:13:43.05" />
                    <SPLIT distance="1300" swimtime="00:14:15.52" />
                    <SPLIT distance="1350" swimtime="00:14:48.39" />
                    <SPLIT distance="1400" swimtime="00:15:21.75" />
                    <SPLIT distance="1450" swimtime="00:15:54.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="507" swimtime="00:02:17.41" resultid="3167" heatid="4753" lane="2" entrytime="00:02:15.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                    <SPLIT distance="150" swimtime="00:01:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="445" swimtime="00:02:18.29" resultid="3168" heatid="4786" lane="2" entrytime="00:02:24.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:07.25" />
                    <SPLIT distance="150" swimtime="00:01:43.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.95" eventid="1971" heatid="4818" lane="3" />
                <ENTRY entrytime="00:04:48.44" eventid="1999" heatid="4861" lane="5" />
                <ENTRY entrytime="00:01:03.32" eventid="2027" heatid="4879" lane="1" />
                <ENTRY entrytime="00:02:11.49" eventid="2041" heatid="4894" lane="5" />
                <ENTRY entrytime="00:04:10.22" eventid="2075" heatid="4911" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Greta Sophie" gender="F" lastname="Westermann" nation="GER" license="274028" athleteid="3174">
              <RESULTS>
                <RESULT eventid="1059" points="552" swimtime="00:01:02.06" resultid="3175" heatid="4670" lane="3" entrytime="00:01:01.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="526" swimtime="00:01:10.20" resultid="3176" heatid="4732" lane="1" entrytime="00:01:12.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="561" swimtime="00:04:44.30" resultid="3177" heatid="4763" lane="1" entrytime="00:04:39.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.28" />
                    <SPLIT distance="150" swimtime="00:01:41.91" />
                    <SPLIT distance="200" swimtime="00:02:18.15" />
                    <SPLIT distance="250" swimtime="00:02:54.78" />
                    <SPLIT distance="300" swimtime="00:03:31.78" />
                    <SPLIT distance="350" swimtime="00:04:08.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="603" swimtime="00:18:08.42" resultid="3178" heatid="4803" lane="2" entrytime="00:18:48.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="150" swimtime="00:01:44.67" />
                    <SPLIT distance="200" swimtime="00:02:21.04" />
                    <SPLIT distance="250" swimtime="00:02:57.70" />
                    <SPLIT distance="300" swimtime="00:03:34.33" />
                    <SPLIT distance="350" swimtime="00:04:10.99" />
                    <SPLIT distance="400" swimtime="00:04:47.98" />
                    <SPLIT distance="450" swimtime="00:05:24.66" />
                    <SPLIT distance="500" swimtime="00:06:01.54" />
                    <SPLIT distance="550" swimtime="00:06:38.18" />
                    <SPLIT distance="600" swimtime="00:07:14.77" />
                    <SPLIT distance="650" swimtime="00:07:51.30" />
                    <SPLIT distance="700" swimtime="00:08:27.83" />
                    <SPLIT distance="750" swimtime="00:09:04.54" />
                    <SPLIT distance="800" swimtime="00:09:40.61" />
                    <SPLIT distance="850" swimtime="00:10:16.83" />
                    <SPLIT distance="900" swimtime="00:10:53.19" />
                    <SPLIT distance="950" swimtime="00:11:29.63" />
                    <SPLIT distance="1000" swimtime="00:12:06.32" />
                    <SPLIT distance="1050" swimtime="00:12:43.22" />
                    <SPLIT distance="1100" swimtime="00:13:19.62" />
                    <SPLIT distance="1150" swimtime="00:13:56.52" />
                    <SPLIT distance="1200" swimtime="00:14:32.32" />
                    <SPLIT distance="1250" swimtime="00:15:08.74" />
                    <SPLIT distance="1300" swimtime="00:15:45.22" />
                    <SPLIT distance="1350" swimtime="00:16:21.49" />
                    <SPLIT distance="1400" swimtime="00:16:57.93" />
                    <SPLIT distance="1450" swimtime="00:17:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1919" points="456" swimtime="00:01:13.58" resultid="5402" heatid="5404" lane="1" entrytime="00:01:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:09:53.98" eventid="2020" heatid="4875" lane="5">
                  <MEETINFO qualificationtime="00:09:53.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.54" eventid="2055" heatid="4904" lane="5" />
                <ENTRY entrytime="00:00:28.32" eventid="2082" heatid="4920" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lea" gender="F" lastname="Winzer" nation="GER" license="316349" athleteid="3182">
              <RESULTS>
                <RESULT eventid="1785" points="433" swimtime="00:01:12.70" resultid="3183" heatid="4719" lane="1" entrytime="00:01:12.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="397" swimtime="00:01:17.08" resultid="3184" heatid="4728" lane="4" entrytime="00:01:15.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="437" swimtime="00:00:32.11" resultid="3185" heatid="4794" lane="4" entrytime="00:00:32.00" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:33.37" eventid="2034" heatid="4885" lane="3" />
                <ENTRY entrytime="00:02:36.02" eventid="2096" heatid="4933" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Simon" gender="M" lastname="Wittner" nation="GER" license="273514" athleteid="3188">
              <RESULTS>
                <RESULT eventid="1820" points="575" swimtime="00:02:11.80" resultid="3189" heatid="4756" lane="5" entrytime="00:02:10.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="100" swimtime="00:01:02.29" />
                    <SPLIT distance="150" swimtime="00:01:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="499" swimtime="00:02:13.09" resultid="3190" heatid="4790" lane="2" entrytime="00:02:11.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                    <SPLIT distance="150" swimtime="00:01:39.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="590" swimtime="00:02:10.70" resultid="5441" heatid="5442" lane="6" entrytime="00:02:11.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                    <SPLIT distance="100" swimtime="00:01:01.42" />
                    <SPLIT distance="150" swimtime="00:01:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="517" swimtime="00:02:11.60" resultid="5497" heatid="4792" lane="6" entrytime="00:02:13.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:04.77" />
                    <SPLIT distance="150" swimtime="00:01:38.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:40.02" eventid="1999" heatid="4862" lane="1" />
                <ENTRY entrytime="00:09:13.63" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:13.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Oliver" gender="M" lastname="Zeidler" nation="GER" license="167736" athleteid="3193">
              <RESULTS>
                <RESULT eventid="1749" points="644" swimtime="00:01:55.02" resultid="3194" heatid="4683" lane="3" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                    <SPLIT distance="100" swimtime="00:00:56.38" />
                    <SPLIT distance="150" swimtime="00:01:26.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="647" swimtime="00:00:23.42" resultid="3195" heatid="4777" lane="5" entrytime="00:00:23.90" />
                <RESULT eventid="1947" points="661" swimtime="00:00:23.25" resultid="5468" heatid="4778" lane="2" entrytime="00:00:23.42" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:50.80" eventid="1971" heatid="4827" lane="3" />
                <ENTRY entrytime="00:01:55.02" eventid="1870" heatid="5342" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="712" swimtime="00:01:41.33" resultid="3197" heatid="4806" lane="3" entrytime="00:01:38.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                    <SPLIT distance="100" swimtime="00:00:53.89" />
                    <SPLIT distance="150" swimtime="00:01:18.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3036" number="1" />
                    <RELAYPOSITION athleteid="3009" number="2" reactiontime="+34" />
                    <RELAYPOSITION athleteid="3072" number="3" reactiontime="+35" />
                    <RELAYPOSITION athleteid="3193" number="4" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:29.29" eventid="2232" heatid="4812" lane="4" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="2062" points="683" swimtime="00:01:58.13" resultid="3199" heatid="4807" lane="3" entrytime="00:01:52.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:02.15" />
                    <SPLIT distance="150" swimtime="00:01:31.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2991" number="1" />
                    <RELAYPOSITION athleteid="3140" number="2" />
                    <RELAYPOSITION athleteid="2972" number="3" />
                    <RELAYPOSITION athleteid="2939" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:42.08" eventid="2224" heatid="4810" lane="3" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6695" nation="GER" region="02" clubid="3452" name="SSG Coburg">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Jonas" gender="M" lastname="Colli" nation="GER" license="257089" athleteid="3453">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.21" eventid="1985" heatid="4844" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Kristof" gender="M" lastname="Kalocsai" nation="GER" license="350499" athleteid="3455">
              <RESULTS>
                <RESULT eventid="1834" points="450" swimtime="00:00:26.43" resultid="3456" heatid="4768" lane="6" entrytime="00:00:26.54" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:59.66" eventid="1971" heatid="4814" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4330" nation="GER" region="02" clubid="2532" name="SSG Neptun Germering e.V.">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Claudia" gender="F" lastname="Dobmeier" nation="GER" license="299888" athleteid="2586">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.85" eventid="2082" heatid="4914" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Mareike" gender="F" lastname="Feller" nation="GER" license="218202" athleteid="2540">
              <RESULTS>
                <RESULT eventid="1785" points="504" swimtime="00:01:09.14" resultid="2541" heatid="4721" lane="2" entrytime="00:01:09.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="488" swimtime="00:01:11.97" resultid="2542" heatid="4733" lane="6" entrytime="00:01:12.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="474" swimtime="00:00:31.25" resultid="2543" heatid="4799" lane="5" entrytime="00:00:30.64" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.20" eventid="2034" heatid="4888" lane="6" />
                <ENTRY entrytime="00:00:28.84" eventid="2082" heatid="4918" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Emily" gender="F" lastname="Gallow" nation="GER" license="384453" athleteid="2593">
              <RESULTS>
                <RESULT eventid="1059" points="500" swimtime="00:01:04.12" resultid="2594" heatid="4663" lane="2" entrytime="00:01:04.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="459" swimtime="00:01:13.45" resultid="2595" heatid="4729" lane="5" entrytime="00:01:14.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="495" swimtime="00:00:30.80" resultid="2596" heatid="4796" lane="4" entrytime="00:00:31.32" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:28.57" eventid="2082" heatid="4919" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Franziska" gender="F" lastname="Godau" nation="GER" license="219095" athleteid="2533">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.37" eventid="2082" heatid="4920" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Miriam" gender="F" lastname="Karcher" nation="GER" license="316822" athleteid="2588">
              <RESULTS>
                <RESULT eventid="1756" points="489" swimtime="00:00:36.54" resultid="2589" heatid="4689" lane="3" entrytime="00:00:36.62" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:22.35" eventid="1992" heatid="4850" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Elisa" gender="F" lastname="Lex" nation="GER" license="323971" athleteid="2591">
              <RESULTS>
                <RESULT eventid="1756" points="459" swimtime="00:00:37.33" resultid="2592" heatid="4688" lane="6" entrytime="00:00:37.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Laura" gender="F" lastname="Obermayer" nation="GER" license="280497" athleteid="2560">
              <RESULTS>
                <RESULT eventid="1756" points="545" swimtime="00:00:35.24" resultid="2561" heatid="4691" lane="2" entrytime="00:00:35.57" />
                <RESULT eventid="1771" points="565" swimtime="00:05:13.79" resultid="2562" heatid="4707" lane="4" entrytime="00:05:16.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:13.11" />
                    <SPLIT distance="150" swimtime="00:01:52.65" />
                    <SPLIT distance="200" swimtime="00:02:34.04" />
                    <SPLIT distance="250" swimtime="00:03:18.20" />
                    <SPLIT distance="300" swimtime="00:04:03.69" />
                    <SPLIT distance="350" swimtime="00:04:39.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="551" swimtime="00:04:46.00" resultid="2563" heatid="4761" lane="3" entrytime="00:04:43.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:07.59" />
                    <SPLIT distance="150" swimtime="00:01:43.71" />
                    <SPLIT distance="200" swimtime="00:02:20.53" />
                    <SPLIT distance="250" swimtime="00:02:57.02" />
                    <SPLIT distance="300" swimtime="00:03:33.79" />
                    <SPLIT distance="350" swimtime="00:04:10.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="492" swimtime="00:02:50.37" resultid="2564" heatid="4783" lane="6" entrytime="00:02:47.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:21.93" />
                    <SPLIT distance="150" swimtime="00:02:06.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:17.49" eventid="1992" heatid="4854" lane="1" />
                <ENTRY entrytime="00:02:27.90" eventid="2055" heatid="4903" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Matthias" gender="M" lastname="Rips" nation="GER" license="226730" athleteid="2546">
              <RESULTS>
                <RESULT eventid="1763" points="538" swimtime="00:01:08.35" resultid="2547" heatid="4697" lane="3" entrytime="00:01:11.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="497" swimtime="00:01:01.15" resultid="2548" heatid="4714" lane="6" entrytime="00:01:00.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="488" swimtime="00:02:19.21" resultid="2549" heatid="4752" lane="4" entrytime="00:02:18.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:47.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.94" eventid="1985" heatid="4846" lane="6" />
                <ENTRY entrytime="00:01:02.64" eventid="2027" heatid="4880" lane="5" />
                <ENTRY entrytime="00:02:29.00" eventid="2089" heatid="4929" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Maximilian" gender="M" lastname="Stadler" nation="GER" license="242037" athleteid="2535">
              <RESULTS>
                <RESULT eventid="1806" points="420" swimtime="00:00:29.66" resultid="2536" heatid="4739" lane="1" entrytime="00:00:30.49" />
                <RESULT eventid="1834" points="432" swimtime="00:00:26.79" resultid="2537" heatid="4766" lane="2" entrytime="00:00:27.32" />
                <RESULT eventid="1848" points="429" swimtime="00:02:19.96" resultid="2538" heatid="4786" lane="4" entrytime="00:02:22.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                    <SPLIT distance="150" swimtime="00:01:42.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:05.68" eventid="2013" heatid="4869" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Nele" gender="F" lastname="Ströbel" nation="GER" license="299265" athleteid="2575">
              <RESULTS>
                <RESULT eventid="1059" points="503" swimtime="00:01:04.00" resultid="2576" heatid="4664" lane="2" entrytime="00:01:03.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="(Zeit: 13:41), Start vor dem Startsignal" eventid="1827" status="DSQ" swimtime="00:04:56.84" resultid="2577" heatid="4759" lane="2" entrytime="00:04:54.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:47.39" />
                    <SPLIT distance="200" swimtime="00:02:25.12" />
                    <SPLIT distance="250" swimtime="00:03:02.55" />
                    <SPLIT distance="300" swimtime="00:03:40.77" />
                    <SPLIT distance="350" swimtime="00:04:19.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="486" swimtime="00:00:31.00" resultid="2578" heatid="4796" lane="6" entrytime="00:00:31.59" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:11.06" eventid="2006" heatid="4863" lane="2" />
                <ENTRY entrytime="00:02:37.51" eventid="2055" heatid="4898" lane="3" />
                <ENTRY entrytime="00:00:29.32" eventid="2082" heatid="4916" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Nikita" gender="M" lastname="Tsvetkov" nation="GER" license="265703" athleteid="2582">
              <RESULTS>
                <RESULT eventid="1806" points="346" swimtime="00:00:31.63" resultid="2583" heatid="4738" lane="2" entrytime="00:00:31.37" />
                <RESULT eventid="1834" points="411" swimtime="00:00:27.23" resultid="2584" heatid="4766" lane="4" entrytime="00:00:27.29" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:59.22" eventid="1971" heatid="4814" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Leopold" gender="M" lastname="Wahl" nation="GER" license="246999" athleteid="2553">
              <RESULTS>
                <RESULT eventid="1778" points="451" swimtime="00:01:03.14" resultid="2554" heatid="4709" lane="3" entrytime="00:01:03.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="447" swimtime="00:00:29.06" resultid="2555" heatid="4742" lane="6" entrytime="00:00:29.13" />
                <RESULT eventid="1848" points="450" swimtime="00:02:17.77" resultid="2556" heatid="4789" lane="2" entrytime="00:02:12.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:07.91" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.94" eventid="1971" heatid="4819" lane="6" />
                <ENTRY entrytime="00:01:02.48" eventid="2013" heatid="4871" lane="6" />
                <ENTRY entrytime="00:00:27.97" eventid="2103" heatid="4942" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Maximilian" gender="M" lastname="Wipplinger" nation="GER" license="293163" athleteid="2567">
              <RESULTS>
                <RESULT eventid="1749" points="601" swimtime="00:01:57.69" resultid="2568" heatid="4682" lane="3" entrytime="00:01:59.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="100" swimtime="00:00:57.30" />
                    <SPLIT distance="150" swimtime="00:01:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1792" points="625" swimtime="00:16:31.56" resultid="2569" heatid="4727" lane="1" entrytime="00:16:36.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="100" swimtime="00:01:01.13" />
                    <SPLIT distance="150" swimtime="00:01:33.36" />
                    <SPLIT distance="200" swimtime="00:02:06.00" />
                    <SPLIT distance="250" swimtime="00:02:39.05" />
                    <SPLIT distance="300" swimtime="00:03:12.29" />
                    <SPLIT distance="350" swimtime="00:03:45.26" />
                    <SPLIT distance="400" swimtime="00:04:18.54" />
                    <SPLIT distance="450" swimtime="00:04:51.98" />
                    <SPLIT distance="500" swimtime="00:05:25.42" />
                    <SPLIT distance="550" swimtime="00:05:58.59" />
                    <SPLIT distance="600" swimtime="00:06:32.08" />
                    <SPLIT distance="650" swimtime="00:07:05.92" />
                    <SPLIT distance="700" swimtime="00:07:39.43" />
                    <SPLIT distance="750" swimtime="00:08:12.75" />
                    <SPLIT distance="800" swimtime="00:08:46.20" />
                    <SPLIT distance="850" swimtime="00:09:19.76" />
                    <SPLIT distance="900" swimtime="00:09:53.50" />
                    <SPLIT distance="950" swimtime="00:10:27.14" />
                    <SPLIT distance="1000" swimtime="00:11:00.28" />
                    <SPLIT distance="1050" swimtime="00:11:33.96" />
                    <SPLIT distance="1100" swimtime="00:12:07.41" />
                    <SPLIT distance="1150" swimtime="00:12:40.75" />
                    <SPLIT distance="1200" swimtime="00:13:14.27" />
                    <SPLIT distance="1250" swimtime="00:13:47.95" />
                    <SPLIT distance="1300" swimtime="00:14:21.21" />
                    <SPLIT distance="1350" swimtime="00:14:54.56" />
                    <SPLIT distance="1400" swimtime="00:15:27.73" />
                    <SPLIT distance="1450" swimtime="00:16:00.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="522" swimtime="00:02:16.12" resultid="2570" heatid="4755" lane="6" entrytime="00:02:12.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:46.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.23" eventid="1971" heatid="4823" lane="3" />
                <ENTRY entrytime="00:04:38.84" eventid="1999" heatid="4862" lane="5" />
                <ENTRY entrytime="00:01:02.71" eventid="2027" heatid="4879" lane="5" />
                <ENTRY entrytime="00:04:09.87" eventid="2075" heatid="4911" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4331" nation="GER" region="02" clubid="3705" name="SSKC Poseidon Aschaffenburg">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Justin" gender="M" lastname="Arapaj" nation="GER" license="243492" swrid="4613309" athleteid="3712">
              <RESULTS>
                <RESULT eventid="1749" points="455" swimtime="00:02:09.17" resultid="3713" heatid="4678" lane="4" entrytime="00:02:06.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="100" swimtime="00:01:00.75" />
                    <SPLIT distance="150" swimtime="00:01:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="467" swimtime="00:02:16.10" resultid="3714" heatid="4787" lane="3" entrytime="00:02:20.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:06.14" />
                    <SPLIT distance="150" swimtime="00:01:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="454" swimtime="00:02:17.40" resultid="5501" heatid="5504" lane="5" entrytime="00:02:16.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                    <SPLIT distance="100" swimtime="00:01:04.54" />
                    <SPLIT distance="150" swimtime="00:01:40.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.73" eventid="1971" heatid="4821" lane="1" />
                <ENTRY entrytime="00:01:04.50" eventid="2013" heatid="4870" lane="1" />
                <ENTRY entrytime="00:00:27.98" eventid="2103" heatid="4942" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Cäcilia" gender="F" lastname="Bausback" nation="GER" license="308503" athleteid="3718">
              <RESULTS>
                <RESULT eventid="1771" points="502" swimtime="00:05:26.28" resultid="3719" heatid="4706" lane="3" entrytime="00:05:29.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                    <SPLIT distance="150" swimtime="00:01:53.41" />
                    <SPLIT distance="200" swimtime="00:02:36.10" />
                    <SPLIT distance="250" swimtime="00:03:23.15" />
                    <SPLIT distance="300" swimtime="00:04:11.56" />
                    <SPLIT distance="350" swimtime="00:04:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="540" swimtime="00:04:47.92" resultid="3720" heatid="4758" lane="4" entrytime="00:04:55.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                    <SPLIT distance="150" swimtime="00:01:43.25" />
                    <SPLIT distance="200" swimtime="00:02:19.74" />
                    <SPLIT distance="250" swimtime="00:02:56.59" />
                    <SPLIT distance="300" swimtime="00:03:34.02" />
                    <SPLIT distance="350" swimtime="00:04:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="458" swimtime="00:00:31.62" resultid="3721" heatid="4793" lane="3" entrytime="00:00:32.11" />
                <RESULT eventid="1905" points="557" swimtime="00:18:37.50" resultid="3722" heatid="4803" lane="5" entrytime="00:18:51.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                    <SPLIT distance="200" swimtime="00:02:21.49" />
                    <SPLIT distance="250" swimtime="00:02:58.59" />
                    <SPLIT distance="300" swimtime="00:03:35.67" />
                    <SPLIT distance="350" swimtime="00:04:13.11" />
                    <SPLIT distance="400" swimtime="00:04:50.43" />
                    <SPLIT distance="450" swimtime="00:05:27.81" />
                    <SPLIT distance="500" swimtime="00:06:05.17" />
                    <SPLIT distance="550" swimtime="00:06:42.65" />
                    <SPLIT distance="600" swimtime="00:07:20.36" />
                    <SPLIT distance="650" swimtime="00:07:57.95" />
                    <SPLIT distance="700" swimtime="00:08:35.80" />
                    <SPLIT distance="750" swimtime="00:09:13.25" />
                    <SPLIT distance="800" swimtime="00:09:51.05" />
                    <SPLIT distance="850" swimtime="00:10:28.75" />
                    <SPLIT distance="900" swimtime="00:11:06.56" />
                    <SPLIT distance="950" swimtime="00:11:44.37" />
                    <SPLIT distance="1000" swimtime="00:12:21.99" />
                    <SPLIT distance="1050" swimtime="00:13:00.11" />
                    <SPLIT distance="1100" swimtime="00:13:37.86" />
                    <SPLIT distance="1150" swimtime="00:14:15.54" />
                    <SPLIT distance="1200" swimtime="00:14:53.17" />
                    <SPLIT distance="1250" swimtime="00:15:30.87" />
                    <SPLIT distance="1300" swimtime="00:16:08.92" />
                    <SPLIT distance="1350" swimtime="00:16:46.57" />
                    <SPLIT distance="1400" swimtime="00:17:24.37" />
                    <SPLIT distance="1450" swimtime="00:18:01.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:10.38" eventid="2006" heatid="4864" lane="5" />
                <ENTRY entrytime="00:02:37.59" eventid="2055" heatid="4898" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Lisa" gender="F" lastname="Diener" nation="GER" license="192721" athleteid="3725">
              <RESULTS>
                <RESULT eventid="1059" points="559" swimtime="00:01:01.77" resultid="3726" heatid="4671" lane="5" entrytime="00:01:01.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="524" swimtime="00:00:30.23" resultid="3727" heatid="4800" lane="5" entrytime="00:00:29.62" />
                <RESULT eventid="1940" points="544" swimtime="00:00:29.85" resultid="5516" heatid="5517" lane="6" entrytime="00:00:30.23" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:28.26" eventid="2082" heatid="4920" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Sebastian" gender="M" lastname="Feser" nation="GER" license="173941" athleteid="3729">
              <RESULTS>
                <RESULT eventid="1778" points="497" swimtime="00:01:01.13" resultid="3730" heatid="4716" lane="6" entrytime="00:01:00.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="399" swimtime="00:00:30.17" resultid="3731" heatid="4740" lane="2" entrytime="00:00:29.34" />
                <RESULT eventid="1834" points="499" swimtime="00:00:25.53" resultid="3732" heatid="4772" lane="4" entrytime="00:00:25.28" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.33" eventid="1971" heatid="4822" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Fabienne" gender="F" lastname="Krüger" nation="GER" license="297473" athleteid="3734">
              <RESULTS>
                <RESULT eventid="1059" points="513" swimtime="00:01:03.58" resultid="3735" heatid="4664" lane="5" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="553" swimtime="00:04:45.66" resultid="3736" heatid="4761" lane="1" entrytime="00:04:48.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:07.52" />
                    <SPLIT distance="150" swimtime="00:01:43.20" />
                    <SPLIT distance="200" swimtime="00:02:19.08" />
                    <SPLIT distance="250" swimtime="00:02:55.55" />
                    <SPLIT distance="300" swimtime="00:03:32.23" />
                    <SPLIT distance="350" swimtime="00:04:09.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:15.75" eventid="1978" heatid="4833" lane="1" />
                <ENTRY entrytime="00:10:14.45" eventid="2020" status="RJC">
                  <MEETINFO qualificationtime="00:10:14.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.42" eventid="2096" heatid="4932" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Dovlat" gender="M" lastname="Mirzoev" nation="GER" license="297743" athleteid="3741">
              <RESULTS>
                <RESULT eventid="1763" points="433" swimtime="00:01:13.48" resultid="3742" heatid="4697" lane="1" entrytime="00:01:13.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="457" swimtime="00:00:26.30" resultid="3743" heatid="4765" lane="2" entrytime="00:00:27.40" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.36" eventid="1971" heatid="4815" lane="2" />
                <ENTRY entrytime="00:00:34.01" eventid="1985" heatid="4841" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Ilyas" gender="M" lastname="Mirzoev" nation="GER" license="297744" athleteid="3746">
              <RESULTS>
                <RESULT eventid="1763" points="386" swimtime="00:01:16.37" resultid="3747" heatid="4696" lane="1" entrytime="00:01:15.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="459" swimtime="00:00:26.26" resultid="3748" heatid="4767" lane="2" entrytime="00:00:26.81" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.80" eventid="1971" heatid="4816" lane="4" />
                <ENTRY entrytime="00:00:28.92" eventid="2103" heatid="4939" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Anna" gender="F" lastname="Reibenspiess" nation="GER" license="297472" athleteid="3751">
              <RESULTS>
                <RESULT eventid="1059" points="616" swimtime="00:00:59.81" resultid="3752" heatid="4673" lane="1" entrytime="00:01:00.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="504" swimtime="00:01:09.11" resultid="3753" heatid="4721" lane="6" entrytime="00:01:10.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="641" swimtime="00:04:31.89" resultid="3754" heatid="4762" lane="3" entrytime="00:04:39.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:39.14" />
                    <SPLIT distance="200" swimtime="00:02:13.57" />
                    <SPLIT distance="250" swimtime="00:02:48.06" />
                    <SPLIT distance="300" swimtime="00:03:23.37" />
                    <SPLIT distance="350" swimtime="00:03:58.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="603" swimtime="00:18:08.47" resultid="3755" heatid="4804" lane="6" entrytime="00:18:21.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                    <SPLIT distance="100" swimtime="00:01:07.66" />
                    <SPLIT distance="150" swimtime="00:01:43.04" />
                    <SPLIT distance="200" swimtime="00:02:18.71" />
                    <SPLIT distance="250" swimtime="00:02:54.07" />
                    <SPLIT distance="300" swimtime="00:03:29.38" />
                    <SPLIT distance="350" swimtime="00:04:05.15" />
                    <SPLIT distance="400" swimtime="00:04:41.14" />
                    <SPLIT distance="450" swimtime="00:05:17.36" />
                    <SPLIT distance="500" swimtime="00:05:53.72" />
                    <SPLIT distance="550" swimtime="00:06:30.18" />
                    <SPLIT distance="600" swimtime="00:07:06.61" />
                    <SPLIT distance="650" swimtime="00:07:43.02" />
                    <SPLIT distance="700" swimtime="00:08:19.58" />
                    <SPLIT distance="750" swimtime="00:08:56.03" />
                    <SPLIT distance="800" swimtime="00:09:32.63" />
                    <SPLIT distance="850" swimtime="00:10:09.62" />
                    <SPLIT distance="900" swimtime="00:10:46.36" />
                    <SPLIT distance="950" swimtime="00:11:23.04" />
                    <SPLIT distance="1000" swimtime="00:11:59.56" />
                    <SPLIT distance="1050" swimtime="00:12:36.62" />
                    <SPLIT distance="1100" swimtime="00:13:13.64" />
                    <SPLIT distance="1150" swimtime="00:13:50.40" />
                    <SPLIT distance="1200" swimtime="00:14:27.58" />
                    <SPLIT distance="1250" swimtime="00:15:04.87" />
                    <SPLIT distance="1300" swimtime="00:15:41.83" />
                    <SPLIT distance="1350" swimtime="00:16:18.75" />
                    <SPLIT distance="1400" swimtime="00:16:55.99" />
                    <SPLIT distance="1450" swimtime="00:17:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="613" swimtime="00:00:59.91" resultid="5326" heatid="5317" lane="2" entrytime="00:00:59.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.48" eventid="1978" heatid="4837" lane="1" />
                <ENTRY entrytime="00:09:35.39" eventid="2020" heatid="4875" lane="4">
                  <MEETINFO qualificationtime="00:09:35.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.86" eventid="2096" heatid="4934" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Niklas" gender="M" lastname="Reibenspiess" nation="GER" license="168669" athleteid="3759">
              <RESULTS>
                <RESULT eventid="1763" points="601" swimtime="00:01:05.86" resultid="3760" heatid="4702" lane="6" entrytime="00:01:06.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="602" swimtime="00:02:09.83" resultid="3761" heatid="4755" lane="1" entrytime="00:02:11.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="100" swimtime="00:01:01.58" />
                    <SPLIT distance="150" swimtime="00:01:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="435" swimtime="00:02:19.32" resultid="3762" heatid="4787" lane="2" entrytime="00:02:21.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                    <SPLIT distance="150" swimtime="00:01:43.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="598" swimtime="00:02:10.11" resultid="5436" heatid="5442" lane="3" entrytime="00:02:09.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                    <SPLIT distance="100" swimtime="00:01:01.73" />
                    <SPLIT distance="150" swimtime="00:01:39.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.08" eventid="1971" heatid="4824" lane="5" />
                <ENTRY entrytime="00:04:47.13" eventid="1999" heatid="4861" lane="2" />
                <ENTRY entrytime="00:02:25.50" eventid="2089" heatid="4928" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Hanna" gender="F" lastname="Seubert" nation="GER" license="257093" athleteid="3766">
              <RESULTS>
                <RESULT eventid="1756" points="503" swimtime="00:00:36.19" resultid="3767" heatid="4692" lane="6" entrytime="00:00:35.43" />
                <RESULT eventid="1785" points="463" swimtime="00:01:11.12" resultid="3768" heatid="4720" lane="5" entrytime="00:01:11.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="449" swimtime="00:02:55.62" resultid="3769" heatid="4780" lane="3" entrytime="00:02:51.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="100" swimtime="00:01:24.86" />
                    <SPLIT distance="150" swimtime="00:02:10.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:18.39" eventid="1992" heatid="4853" lane="4" />
                <ENTRY entrytime="00:00:33.42" eventid="2034" heatid="4885" lane="2" />
                <ENTRY entrytime="00:00:28.10" eventid="2082" heatid="4921" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Philipp" gender="M" lastname="Walter" nation="GER" license="284784" athleteid="3773">
              <RESULTS>
                <RESULT eventid="1749" points="506" swimtime="00:02:04.62" resultid="3774" heatid="4678" lane="6" entrytime="00:02:07.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="100" swimtime="00:01:00.00" />
                    <SPLIT distance="150" swimtime="00:01:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1792" points="511" swimtime="00:17:40.14" resultid="3775" heatid="4726" lane="5" entrytime="00:17:51.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:03.94" />
                    <SPLIT distance="150" swimtime="00:01:38.47" />
                    <SPLIT distance="200" swimtime="00:02:13.54" />
                    <SPLIT distance="250" swimtime="00:02:48.61" />
                    <SPLIT distance="300" swimtime="00:03:24.08" />
                    <SPLIT distance="350" swimtime="00:03:59.74" />
                    <SPLIT distance="400" swimtime="00:04:34.85" />
                    <SPLIT distance="450" swimtime="00:05:10.33" />
                    <SPLIT distance="500" swimtime="00:05:46.17" />
                    <SPLIT distance="550" swimtime="00:06:21.70" />
                    <SPLIT distance="600" swimtime="00:06:57.23" />
                    <SPLIT distance="650" swimtime="00:07:32.86" />
                    <SPLIT distance="700" swimtime="00:08:08.41" />
                    <SPLIT distance="750" swimtime="00:08:44.35" />
                    <SPLIT distance="800" swimtime="00:09:20.22" />
                    <SPLIT distance="850" swimtime="00:09:56.28" />
                    <SPLIT distance="900" swimtime="00:10:32.31" />
                    <SPLIT distance="950" swimtime="00:11:08.51" />
                    <SPLIT distance="1000" swimtime="00:11:44.57" />
                    <SPLIT distance="1050" swimtime="00:12:20.84" />
                    <SPLIT distance="1100" swimtime="00:12:56.85" />
                    <SPLIT distance="1150" swimtime="00:13:32.66" />
                    <SPLIT distance="1200" swimtime="00:14:08.78" />
                    <SPLIT distance="1250" swimtime="00:14:44.44" />
                    <SPLIT distance="1300" swimtime="00:15:19.89" />
                    <SPLIT distance="1350" swimtime="00:15:55.67" />
                    <SPLIT distance="1400" swimtime="00:16:31.47" />
                    <SPLIT distance="1450" swimtime="00:17:06.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="395" swimtime="00:00:30.27" resultid="3776" heatid="4739" lane="6" entrytime="00:00:30.72" />
                <RESULT eventid="1848" points="445" swimtime="00:02:18.26" resultid="3777" heatid="4788" lane="5" entrytime="00:02:18.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:06.31" />
                    <SPLIT distance="150" swimtime="00:01:42.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:58.00" eventid="1999" heatid="4860" lane="3" />
                <ENTRY entrytime="00:04:31.31" eventid="2075" heatid="4908" lane="4" />
                <ENTRY entrytime="00:09:16.88" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:16.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="508" swimtime="00:01:53.41" resultid="3781" heatid="4805" lane="2" entrytime="00:01:54.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:28.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3729" number="1" />
                    <RELAYPOSITION athleteid="3759" number="2" reactiontime="+44" />
                    <RELAYPOSITION athleteid="3746" number="3" reactiontime="+38" />
                    <RELAYPOSITION athleteid="3712" number="4" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:42.43" eventid="2232" heatid="4811" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3729" number="1" />
                    <RELAYPOSITION athleteid="3759" number="2" />
                    <RELAYPOSITION athleteid="3712" number="3" />
                    <RELAYPOSITION athleteid="3746" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="2062" points="540" swimtime="00:02:07.69" resultid="3783" heatid="4807" lane="6" entrytime="00:02:10.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3751" number="1" />
                    <RELAYPOSITION athleteid="3766" number="2" />
                    <RELAYPOSITION athleteid="3718" number="3" />
                    <RELAYPOSITION athleteid="3725" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:55.78" eventid="2224" heatid="4810" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3725" number="1" />
                    <RELAYPOSITION athleteid="3751" number="2" />
                    <RELAYPOSITION athleteid="3766" number="3" />
                    <RELAYPOSITION athleteid="3734" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4347" nation="GER" region="02" clubid="4572" name="SV Bayreuth">
          <ATHLETES>
            <ATHLETE birthdate="1991-01-01" firstname="Christoph" gender="M" lastname="Argauer" nation="GER" license="134500" athleteid="4573">
              <RESULTS>
                <RESULT eventid="1749" points="465" swimtime="00:02:08.23" resultid="4574" heatid="4680" lane="2" entrytime="00:02:03.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="100" swimtime="00:00:59.81" />
                    <SPLIT distance="150" swimtime="00:01:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1763" points="448" swimtime="00:01:12.67" resultid="4575" heatid="4699" lane="3" entrytime="00:01:09.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.32" eventid="1971" heatid="4820" lane="4" />
                <ENTRY entrytime="00:00:32.10" eventid="1985" heatid="4844" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Jette" gender="F" lastname="Barthmann" nation="GER" license="297427" athleteid="4578">
              <RESULTS>
                <RESULT eventid="1785" points="408" swimtime="00:01:14.15" resultid="4579" heatid="4719" lane="6" entrytime="00:01:13.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="471" swimtime="00:00:31.32" resultid="4580" heatid="4796" lane="3" entrytime="00:00:31.21" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:10.73" eventid="2006" heatid="4863" lane="3" />
                <ENTRY entrytime="00:00:34.09" eventid="2034" heatid="4884" lane="6" />
                <ENTRY entrytime="00:02:37.31" eventid="2055" heatid="4899" lane="6" />
                <ENTRY entrytime="00:02:36.81" eventid="2096" heatid="4932" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Marc Oliver" gender="M" lastname="Birkle" nation="GER" license="269134" athleteid="4585">
              <RESULTS>
                <RESULT eventid="1749" points="483" swimtime="00:02:06.58" resultid="4586" heatid="4678" lane="3" entrytime="00:02:05.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="100" swimtime="00:00:59.60" />
                    <SPLIT distance="150" swimtime="00:01:32.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="451" swimtime="00:00:26.41" resultid="4587" heatid="4769" lane="3" entrytime="00:00:26.05" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.95" eventid="1971" heatid="4818" lane="4" />
                <ENTRY entrytime="00:00:32.78" eventid="1985" heatid="4842" lane="3" />
                <ENTRY entrytime="00:04:33.07" eventid="2075" heatid="4908" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Maximilian" gender="M" lastname="Deichsel" nation="GER" license="138788" athleteid="4591">
              <RESULTS>
                <RESULT eventid="1778" points="549" swimtime="00:00:59.14" resultid="4592" heatid="4715" lane="6" entrytime="00:01:00.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="590" swimtime="00:02:10.71" resultid="4593" heatid="4754" lane="5" entrytime="00:02:11.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                    <SPLIT distance="100" swimtime="00:01:01.48" />
                    <SPLIT distance="150" swimtime="00:01:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5369" points="553" swimtime="00:00:59.00" resultid="5376" heatid="5378" lane="3" entrytime="00:00:59.14" />
                <RESULT eventid="1926" points="577" swimtime="00:02:11.62" resultid="5437" heatid="5442" lane="4" entrytime="00:02:10.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:01:01.48" />
                    <SPLIT distance="150" swimtime="00:01:40.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:45.15" eventid="1999" heatid="4861" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Carmen" gender="F" lastname="Gräbner" nation="GER" license="297780" athleteid="4595">
              <RESULTS>
                <RESULT eventid="1756" points="468" swimtime="00:00:37.08" resultid="4596" heatid="4689" lane="2" entrytime="00:00:36.85" />
                <RESULT eventid="1771" points="476" swimtime="00:05:32.28" resultid="4597" heatid="4707" lane="5" entrytime="00:05:27.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:02:00.69" />
                    <SPLIT distance="200" swimtime="00:02:45.87" />
                    <SPLIT distance="250" swimtime="00:03:29.98" />
                    <SPLIT distance="300" swimtime="00:04:17.27" />
                    <SPLIT distance="350" swimtime="00:04:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="464" swimtime="00:02:53.74" resultid="4598" heatid="4781" lane="1" entrytime="00:02:50.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:01:23.48" />
                    <SPLIT distance="150" swimtime="00:02:09.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:19.50" eventid="1992" heatid="4852" lane="5" />
                <ENTRY entrytime="00:02:33.85" eventid="2055" heatid="4901" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Nico" gender="M" lastname="Heilmann" nation="GER" license="291040" athleteid="4601">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.72" eventid="1985" heatid="4840" lane="3" />
                <ENTRY entrytime="00:02:42.39" eventid="2089" heatid="4925" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Luisa" gender="F" lastname="Kauper" nation="GER" license="305148" athleteid="4604">
              <RESULTS>
                <RESULT eventid="1756" points="494" swimtime="00:00:36.41" resultid="4605" heatid="4687" lane="2" entrytime="00:00:37.71" />
                <RESULT eventid="1841" points="513" swimtime="00:02:48.08" resultid="4606" heatid="4781" lane="3" entrytime="00:02:48.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:21.49" />
                    <SPLIT distance="150" swimtime="00:02:05.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:20.46" eventid="1992" heatid="4851" lane="2" />
                <ENTRY entrytime="00:02:35.98" eventid="2055" heatid="4899" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Florian" gender="M" lastname="Müller" nation="GER" license="266235" athleteid="4609">
              <RESULTS>
                <RESULT eventid="1763" points="566" swimtime="00:01:07.22" resultid="4610" heatid="4703" lane="6" entrytime="00:01:06.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="490" swimtime="00:01:01.41" resultid="4611" heatid="4713" lane="3" entrytime="00:01:00.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="541" swimtime="00:02:14.50" resultid="4612" heatid="4753" lane="3" entrytime="00:02:14.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                    <SPLIT distance="100" swimtime="00:01:05.98" />
                    <SPLIT distance="150" swimtime="00:01:43.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.14" eventid="1971" heatid="4822" lane="4" />
                <ENTRY entrytime="00:00:31.16" eventid="1985" heatid="4845" lane="1" />
                <ENTRY entrytime="00:02:23.81" eventid="2089" heatid="4929" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Selina" gender="F" lastname="Müller" nation="GER" license="242742" athleteid="4616">
              <RESULTS>
                <RESULT eventid="1785" points="482" swimtime="00:01:10.18" resultid="4617" heatid="4724" lane="6" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.77" eventid="2034" heatid="4888" lane="1" />
                <ENTRY entrytime="00:02:24.16" eventid="2096" heatid="4936" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Stefanie" gender="F" lastname="Raps" nation="GER" license="234205" athleteid="4620">
              <RESULTS>
                <RESULT eventid="1813" points="503" swimtime="00:02:30.37" resultid="4621" heatid="4746" lane="1" entrytime="00:02:34.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                    <SPLIT distance="150" swimtime="00:01:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="522" swimtime="00:04:51.22" resultid="4622" heatid="4760" lane="6" entrytime="00:04:52.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:47.12" />
                    <SPLIT distance="200" swimtime="00:02:24.28" />
                    <SPLIT distance="250" swimtime="00:03:01.50" />
                    <SPLIT distance="300" swimtime="00:03:38.78" />
                    <SPLIT distance="350" swimtime="00:04:16.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1933" points="521" swimtime="00:02:28.60" resultid="5427" heatid="5429" lane="5" entrytime="00:02:30.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                    <SPLIT distance="150" swimtime="00:01:50.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:21.48" eventid="1978" heatid="4829" lane="5" />
                <ENTRY entrytime="00:01:11.67" eventid="2006" heatid="4863" lane="5" />
                <ENTRY entrytime="00:02:34.79" eventid="2055" heatid="4900" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="515" swimtime="00:01:52.85" resultid="4626" heatid="4805" lane="4" entrytime="00:01:54.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="100" swimtime="00:01:01.14" />
                    <SPLIT distance="150" swimtime="00:01:27.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4591" number="1" />
                    <RELAYPOSITION athleteid="4573" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="4609" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="4585" number="4" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:44.00" eventid="2232" heatid="4811" lane="2" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4356" nation="GER" region="02" clubid="2436" name="SV GR.-W. Holzkirchen">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-01" firstname="Ludwig" gender="M" lastname="Huber" nation="GER" license="181978" athleteid="2437">
              <RESULTS>
                <RESULT eventid="1749" points="555" swimtime="00:02:00.87" resultid="2438" heatid="4682" lane="6" entrytime="00:02:01.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                    <SPLIT distance="100" swimtime="00:00:56.99" />
                    <SPLIT distance="150" swimtime="00:01:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1763" points="441" swimtime="00:01:13.05" resultid="2439" heatid="4698" lane="4" entrytime="00:01:10.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="506" swimtime="00:01:00.76" resultid="2440" heatid="4713" lane="6" entrytime="00:01:01.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="582" swimtime="00:00:24.26" resultid="2441" heatid="4776" lane="6" entrytime="00:00:24.54" />
                <RESULT eventid="5443" points="567" swimtime="00:00:24.47" resultid="5451" heatid="5452" lane="4" entrytime="00:00:24.26" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.20" eventid="1971" heatid="4824" lane="6" />
                <ENTRY entrytime="00:00:32.00" eventid="1985" heatid="4844" lane="5" />
                <ENTRY entrytime="00:00:27.26" eventid="2103" heatid="4944" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5713" nation="GER" region="02" clubid="2488" name="SV Hengersberg">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Fabian" gender="M" lastname="Miller" nation="GER" license="282389" athleteid="2489">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.08" eventid="1971" heatid="4815" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Erik" gender="M" lastname="Stögbauer" nation="GER" license="291450" athleteid="2491">
              <RESULTS>
                <RESULT eventid="1806" points="369" swimtime="00:00:30.97" resultid="2492" heatid="4738" lane="4" entrytime="00:00:31.16" />
                <RESULT eventid="1834" points="429" swimtime="00:00:26.86" resultid="2493" heatid="4767" lane="6" entrytime="00:00:27.00" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:00.13" eventid="1971" heatid="4813" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4341" nation="GER" region="02" clubid="4628" name="SV Hof 1911 e. V.">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Leon" gender="M" lastname="Richter" nation="GER" license="270159" athleteid="4636">
              <RESULTS>
                <RESULT eventid="1792" points="436" swimtime="00:18:37.95" resultid="4637" heatid="4726" lane="1" entrytime="00:18:47.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                    <SPLIT distance="100" swimtime="00:01:04.65" />
                    <SPLIT distance="150" swimtime="00:01:41.42" />
                    <SPLIT distance="200" swimtime="00:02:18.94" />
                    <SPLIT distance="250" swimtime="00:02:55.96" />
                    <SPLIT distance="300" swimtime="00:03:33.62" />
                    <SPLIT distance="350" swimtime="00:04:11.68" />
                    <SPLIT distance="400" swimtime="00:04:49.72" />
                    <SPLIT distance="450" swimtime="00:05:27.00" />
                    <SPLIT distance="500" swimtime="00:06:04.96" />
                    <SPLIT distance="550" swimtime="00:06:42.30" />
                    <SPLIT distance="600" swimtime="00:07:20.25" />
                    <SPLIT distance="650" swimtime="00:07:57.96" />
                    <SPLIT distance="700" swimtime="00:08:35.73" />
                    <SPLIT distance="750" swimtime="00:09:14.02" />
                    <SPLIT distance="800" swimtime="00:09:51.78" />
                    <SPLIT distance="850" swimtime="00:10:30.58" />
                    <SPLIT distance="900" swimtime="00:11:08.48" />
                    <SPLIT distance="950" swimtime="00:11:45.99" />
                    <SPLIT distance="1000" swimtime="00:12:24.48" />
                    <SPLIT distance="1050" swimtime="00:13:02.65" />
                    <SPLIT distance="1100" swimtime="00:13:40.91" />
                    <SPLIT distance="1150" swimtime="00:14:18.61" />
                    <SPLIT distance="1200" swimtime="00:14:56.60" />
                    <SPLIT distance="1250" swimtime="00:15:35.03" />
                    <SPLIT distance="1300" swimtime="00:16:12.39" />
                    <SPLIT distance="1350" swimtime="00:16:50.58" />
                    <SPLIT distance="1400" swimtime="00:17:27.84" />
                    <SPLIT distance="1450" swimtime="00:18:04.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="430" swimtime="00:00:26.83" resultid="4638" heatid="4767" lane="1" entrytime="00:00:26.95" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:59.88" eventid="1971" heatid="4814" lane="6" />
                <ENTRY entrytime="00:04:39.47" eventid="2075" heatid="4906" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Matthias" gender="M" lastname="Schmidt" nation="GER" license="209569" athleteid="4641">
              <RESULTS>
                <RESULT eventid="1834" points="443" swimtime="00:00:26.56" resultid="4642" heatid="4768" lane="4" entrytime="00:00:26.33" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:27.80" eventid="2103" heatid="4942" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4364" nation="GER" region="02" clubid="3247" name="SV Ottobrunn 1970 e.V.">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Birte" gender="F" lastname="Schiemann" nation="GER" license="260141" athleteid="3248">
              <ENTRIES>
                <ENTRY entrytime="00:02:19.40" eventid="1978" heatid="4831" lane="5" />
                <ENTRY entrytime="00:00:33.00" eventid="2034" heatid="4886" lane="6" />
                <ENTRY entrytime="00:00:28.76" eventid="2082" heatid="4918" lane="2" />
                <ENTRY entrytime="00:02:32.49" eventid="2096" heatid="4934" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4384" nation="GER" region="02" clubid="2445" name="SV Wacker Burghausen">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Verena" gender="F" lastname="Bergmann" nation="GER" license="295270" athleteid="2446">
              <RESULTS>
                <RESULT eventid="1785" points="438" swimtime="00:01:12.46" resultid="2447" heatid="4719" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="450" swimtime="00:01:13.91" resultid="2448" heatid="4730" lane="3" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Yannick" gender="M" lastname="Buschhardt" nation="GER" license="227101" athleteid="2449">
              <RESULTS>
                <RESULT eventid="1806" points="538" swimtime="00:00:27.31" resultid="2450" heatid="4742" lane="2" entrytime="00:00:28.00" />
                <RESULT eventid="1834" points="555" swimtime="00:00:24.64" resultid="2451" heatid="4777" lane="6" entrytime="00:00:24.50" />
                <RESULT eventid="1912" points="532" swimtime="00:00:27.41" resultid="5407" heatid="4744" lane="2" entrytime="00:00:27.31" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.60" eventid="1971" heatid="4825" lane="6" />
                <ENTRY entrytime="00:00:59.00" eventid="2013" heatid="4872" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Marina" gender="F" lastname="Hammerl" nation="GER" license="284445" athleteid="2454">
              <RESULTS>
                <RESULT eventid="1059" points="554" swimtime="00:01:01.95" resultid="2455" heatid="4668" lane="5" entrytime="00:01:02.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1813" points="510" swimtime="00:02:29.62" resultid="2456" heatid="4747" lane="1" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="519" swimtime="00:00:30.33" resultid="2457" heatid="4797" lane="3" entrytime="00:00:31.00" />
                <RESULT eventid="1933" points="511" swimtime="00:02:29.53" resultid="5425" heatid="5429" lane="4" entrytime="00:02:29.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:10.77" />
                    <SPLIT distance="150" swimtime="00:01:51.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:16.50" eventid="1978" heatid="4832" lane="4" />
                <ENTRY entrytime="00:01:08.00" eventid="2006" heatid="4867" lane="6" />
                <ENTRY entrytime="00:00:29.50" eventid="2082" heatid="4915" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Dominik" gender="M" lastname="Kohlschmid" nation="GER" license="242746" athleteid="2461">
              <RESULTS>
                <RESULT eventid="1763" points="598" swimtime="00:01:05.98" resultid="2462" heatid="4701" lane="5" entrytime="00:01:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="581" swimtime="00:00:58.05" resultid="2463" heatid="4716" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="628" swimtime="00:02:08.00" resultid="2464" heatid="4754" lane="4" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="100" swimtime="00:01:01.03" />
                    <SPLIT distance="150" swimtime="00:01:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="594" swimtime="00:02:10.36" resultid="5435" heatid="4757" lane="6" entrytime="00:02:08.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1898" points="619" swimtime="00:00:56.82" resultid="5457" heatid="4717" lane="1" entrytime="00:00:58.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.40" eventid="1971" heatid="4823" lane="2" />
                <ENTRY entrytime="00:00:30.00" eventid="1985" heatid="4846" lane="5" />
                <ENTRY entrytime="00:00:59.00" eventid="2027" heatid="4880" lane="4" />
                <ENTRY entrytime="00:02:27.00" eventid="2089" heatid="4928" lane="1" />
                <ENTRY entrytime="00:00:27.00" eventid="2103" heatid="4947" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Paulina" gender="F" lastname="Sandner" nation="GER" license="316586" athleteid="2470">
              <RESULTS>
                <RESULT eventid="1059" points="566" swimtime="00:01:01.51" resultid="2471" heatid="4668" lane="4" entrytime="00:01:02.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="513" swimtime="00:00:35.96" resultid="2472" heatid="4691" lane="1" entrytime="00:00:35.70" />
                <RESULT eventid="1799" points="528" swimtime="00:01:10.08" resultid="2473" heatid="4735" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1919" points="536" swimtime="00:01:09.76" resultid="5401" heatid="5404" lane="5" entrytime="00:01:10.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:17.00" eventid="1992" heatid="4854" lane="3" />
                <ENTRY entrytime="00:00:29.00" eventid="2082" heatid="4917" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Marlene" gender="F" lastname="Sommoggy von" nation="GER" license="304160" athleteid="2476">
              <RESULTS>
                <RESULT eventid="1756" points="598" swimtime="00:00:34.18" resultid="2477" heatid="4690" lane="3" entrytime="00:00:36.00" />
                <RESULT eventid="1799" points="490" swimtime="00:01:11.88" resultid="2478" heatid="4733" lane="2" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="549" swimtime="00:02:44.28" resultid="2479" heatid="4782" lane="6" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:19.76" />
                    <SPLIT distance="150" swimtime="00:02:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1877" points="592" swimtime="00:00:34.29" resultid="5351" heatid="5355" lane="2" entrytime="00:00:34.18" />
                <RESULT eventid="1954" points="562" swimtime="00:02:43.04" resultid="5489" heatid="5491" lane="1" entrytime="00:02:44.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="150" swimtime="00:02:02.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:17.00" eventid="1992" heatid="4854" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4387" nation="GER" region="02" clubid="4648" name="SV Weiden">
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Lisa" gender="F" lastname="Biersack" nation="GER" license="225273" athleteid="4649">
              <RESULTS>
                <RESULT eventid="1785" points="553" swimtime="00:01:07.04" resultid="4650" heatid="4724" lane="4" entrytime="00:01:04.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="470" swimtime="00:01:12.85" resultid="4651" heatid="4736" lane="1" entrytime="00:01:10.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="485" swimtime="00:00:31.03" resultid="4652" heatid="4800" lane="6" entrytime="00:00:29.92" />
                <RESULT eventid="1891" points="534" swimtime="00:01:07.80" resultid="5389" heatid="5391" lane="1" entrytime="00:01:07.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.02" eventid="2034" heatid="4887" lane="2" />
                <ENTRY entrytime="00:02:23.95" eventid="2096" heatid="4935" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Alina" gender="F" lastname="Zimmermann" nation="GER" license="193325" athleteid="4655">
              <RESULTS>
                <RESULT eventid="1059" points="537" swimtime="00:01:02.62" resultid="4656" heatid="4671" lane="4" entrytime="00:01:01.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="458" swimtime="00:01:13.51" resultid="4657" heatid="4734" lane="6" entrytime="00:01:11.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="467" swimtime="00:00:31.41" resultid="4658" heatid="4799" lane="3" entrytime="00:00:30.49" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:12.72" eventid="1978" heatid="4835" lane="5" />
                <ENTRY entrytime="00:01:07.53" eventid="2006" heatid="4866" lane="1" />
                <ENTRY entrytime="00:00:28.03" eventid="2082" heatid="4923" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4339" nation="GER" region="02" clubid="3493" name="SV Würzburg 05">
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Leonie Antonia" gender="F" lastname="Beck" nation="GER" license="186145" athleteid="3502">
              <RESULTS>
                <RESULT eventid="1059" points="695" swimtime="00:00:57.46" resultid="3503" heatid="4674" lane="3" entrytime="00:00:55.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="679" swimtime="00:02:33.07" resultid="3504" heatid="4784" lane="3" entrytime="00:02:27.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="719" swimtime="00:00:56.82" resultid="5318" heatid="4675" lane="3" entrytime="00:00:57.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1954" points="732" swimtime="00:02:29.26" resultid="5479" heatid="4785" lane="3" entrytime="00:02:33.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:57.90" eventid="1978" heatid="4838" lane="3" />
                <ENTRY entrytime="00:02:11.87" eventid="2055" heatid="4904" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Maximilian" gender="M" lastname="Beck" nation="GER" license="161820" athleteid="3507">
              <RESULTS>
                <RESULT eventid="1763" points="650" swimtime="00:01:04.19" resultid="3508" heatid="4702" lane="3" entrytime="00:01:02.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="650" swimtime="00:02:06.51" resultid="3509" heatid="4756" lane="3" entrytime="00:02:03.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="100" swimtime="00:01:01.52" />
                    <SPLIT distance="150" swimtime="00:01:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="583" swimtime="00:00:24.24" resultid="3510" heatid="4775" lane="2" entrytime="00:00:23.65" />
                <RESULT eventid="1884" points="660" swimtime="00:01:03.86" resultid="5361" heatid="4704" lane="6" entrytime="00:01:04.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="650" swimtime="00:02:06.51" resultid="5431" heatid="4757" lane="4" entrytime="00:02:06.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="100" swimtime="00:01:01.58" />
                    <SPLIT distance="150" swimtime="00:01:37.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.13" eventid="1985" heatid="4847" lane="4" />
                <ENTRY entrytime="00:00:57.94" eventid="2027" heatid="4880" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Sebastian Aurelius" gender="M" lastname="Beck" nation="GER" license="236295" athleteid="3513">
              <RESULTS>
                <RESULT eventid="1749" points="646" swimtime="00:01:54.95" resultid="3514" heatid="4683" lane="4" entrytime="00:01:53.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.71" />
                    <SPLIT distance="100" swimtime="00:00:56.38" />
                    <SPLIT distance="150" swimtime="00:01:26.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="633" swimtime="00:02:07.63" resultid="3515" heatid="4755" lane="4" entrytime="00:02:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="100" swimtime="00:01:00.88" />
                    <SPLIT distance="150" swimtime="00:01:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="653" swimtime="00:02:06.36" resultid="5433" heatid="4757" lane="5" entrytime="00:02:07.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                    <SPLIT distance="150" swimtime="00:01:38.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:52.39" eventid="1971" heatid="4825" lane="2" />
                <ENTRY entrytime="00:03:58.67" eventid="2075" heatid="4912" lane="2" />
                <ENTRY entrytime="00:08:30.03" eventid="2168" heatid="4809" lane="1">
                  <MEETINFO qualificationtime="00:08:30.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.95" eventid="1870" heatid="5342" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Max" gender="M" lastname="Brandenstein" nation="GER" license="312913" athleteid="3519">
              <RESULTS>
                <RESULT eventid="1792" points="605" swimtime="00:16:42.40" resultid="3520" heatid="4727" lane="6" entrytime="00:16:41.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:01.13" />
                    <SPLIT distance="150" swimtime="00:01:33.85" />
                    <SPLIT distance="200" swimtime="00:02:06.76" />
                    <SPLIT distance="250" swimtime="00:02:39.78" />
                    <SPLIT distance="300" swimtime="00:03:13.01" />
                    <SPLIT distance="350" swimtime="00:03:46.47" />
                    <SPLIT distance="400" swimtime="00:04:20.02" />
                    <SPLIT distance="450" swimtime="00:04:53.51" />
                    <SPLIT distance="500" swimtime="00:05:27.08" />
                    <SPLIT distance="550" swimtime="00:06:00.59" />
                    <SPLIT distance="600" swimtime="00:06:34.58" />
                    <SPLIT distance="650" swimtime="00:07:08.47" />
                    <SPLIT distance="700" swimtime="00:07:42.14" />
                    <SPLIT distance="750" swimtime="00:08:16.03" />
                    <SPLIT distance="800" swimtime="00:08:49.85" />
                    <SPLIT distance="850" swimtime="00:09:23.59" />
                    <SPLIT distance="900" swimtime="00:09:57.78" />
                    <SPLIT distance="950" swimtime="00:10:31.62" />
                    <SPLIT distance="1000" swimtime="00:11:05.55" />
                    <SPLIT distance="1050" swimtime="00:11:39.29" />
                    <SPLIT distance="1100" swimtime="00:12:13.22" />
                    <SPLIT distance="1150" swimtime="00:12:47.11" />
                    <SPLIT distance="1200" swimtime="00:13:20.90" />
                    <SPLIT distance="1250" swimtime="00:13:54.84" />
                    <SPLIT distance="1300" swimtime="00:14:28.99" />
                    <SPLIT distance="1350" swimtime="00:15:02.75" />
                    <SPLIT distance="1400" swimtime="00:15:36.48" />
                    <SPLIT distance="1450" swimtime="00:16:09.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="449" swimtime="00:00:26.45" resultid="3521" heatid="4769" lane="6" entrytime="00:00:26.30" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.74" eventid="1971" heatid="4819" lane="4" />
                <ENTRY entrytime="00:04:11.51" eventid="2075" heatid="4910" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Frederik" gender="M" lastname="Bär" nation="GER" license="249941" athleteid="3497">
              <RESULTS>
                <RESULT eventid="1806" points="512" swimtime="00:00:27.77" resultid="3498" heatid="4741" lane="5" entrytime="00:00:28.50" />
                <RESULT eventid="1834" points="557" swimtime="00:00:24.62" resultid="3499" heatid="4774" lane="2" entrytime="00:00:24.78" />
                <RESULT eventid="1912" points="509" swimtime="00:00:27.82" resultid="5412" heatid="5417" lane="4" entrytime="00:00:27.77" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="1971" heatid="4823" lane="6" />
                <ENTRY entrytime="00:01:02.00" eventid="2027" heatid="4881" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Klemens" gender="M" lastname="Degenhardt" nation="GER" license="140643" athleteid="3524">
              <RESULTS>
                <RESULT eventid="1763" points="656" swimtime="00:01:03.99" resultid="3525" heatid="4703" lane="3" entrytime="00:01:00.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="523" swimtime="00:02:11.10" resultid="3526" heatid="4791" lane="1" entrytime="00:02:14.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:04.17" />
                    <SPLIT distance="150" swimtime="00:01:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1884" points="670" swimtime="00:01:03.54" resultid="5359" heatid="4704" lane="5" entrytime="00:01:03.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:28.04" eventid="1985" heatid="4847" lane="3" />
                <ENTRY entrytime="00:02:12.26" eventid="2089" heatid="4930" lane="3" />
                <ENTRY entrytime="00:08:34.84" eventid="2168" heatid="4808" lane="3">
                  <MEETINFO qualificationtime="00:08:34.84" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Carolin" gender="F" lastname="Dorfner" nation="GER" license="244045" athleteid="3530">
              <RESULTS>
                <RESULT eventid="1059" points="626" swimtime="00:00:59.51" resultid="3531" heatid="4673" lane="2" entrytime="00:00:59.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1813" points="647" swimtime="00:02:18.28" resultid="3532" heatid="4746" lane="4" entrytime="00:02:19.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="597" swimtime="00:00:28.94" resultid="3533" heatid="4801" lane="5" entrytime="00:00:29.55" />
                <RESULT eventid="1863" points="621" swimtime="00:00:59.65" resultid="5324" heatid="5317" lane="3" entrytime="00:00:59.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1933" points="649" swimtime="00:02:18.13" resultid="5418" heatid="4748" lane="3" entrytime="00:02:18.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                    <SPLIT distance="100" swimtime="00:01:06.58" />
                    <SPLIT distance="150" swimtime="00:01:42.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:03.53" eventid="2006" heatid="4867" lane="4" />
                <ENTRY entrytime="00:02:21.52" eventid="2055" heatid="4904" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Romy" gender="F" lastname="Dreher" nation="GER" license="269748" athleteid="3546">
              <RESULTS>
                <RESULT eventid="1059" points="603" swimtime="00:01:00.24" resultid="3547" heatid="4672" lane="5" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="650" swimtime="00:04:30.70" resultid="3548" heatid="4764" lane="2" entrytime="00:04:22.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:01:04.62" />
                    <SPLIT distance="150" swimtime="00:01:38.82" />
                    <SPLIT distance="200" swimtime="00:02:12.99" />
                    <SPLIT distance="250" swimtime="00:02:47.00" />
                    <SPLIT distance="300" swimtime="00:03:21.62" />
                    <SPLIT distance="350" swimtime="00:03:56.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="686" swimtime="00:17:22.76" resultid="3549" heatid="4804" lane="2" entrytime="00:17:40.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                    <SPLIT distance="150" swimtime="00:01:41.56" />
                    <SPLIT distance="200" swimtime="00:02:16.32" />
                    <SPLIT distance="250" swimtime="00:02:51.27" />
                    <SPLIT distance="300" swimtime="00:03:26.17" />
                    <SPLIT distance="350" swimtime="00:04:01.29" />
                    <SPLIT distance="400" swimtime="00:04:36.47" />
                    <SPLIT distance="450" swimtime="00:05:11.57" />
                    <SPLIT distance="500" swimtime="00:05:46.66" />
                    <SPLIT distance="550" swimtime="00:06:21.45" />
                    <SPLIT distance="600" swimtime="00:06:56.25" />
                    <SPLIT distance="650" swimtime="00:07:31.16" />
                    <SPLIT distance="700" swimtime="00:08:06.36" />
                    <SPLIT distance="750" swimtime="00:08:41.27" />
                    <SPLIT distance="800" swimtime="00:09:16.34" />
                    <SPLIT distance="850" swimtime="00:09:51.19" />
                    <SPLIT distance="900" swimtime="00:10:26.30" />
                    <SPLIT distance="950" swimtime="00:11:01.19" />
                    <SPLIT distance="1000" swimtime="00:11:36.39" />
                    <SPLIT distance="1050" swimtime="00:12:11.37" />
                    <SPLIT distance="1100" swimtime="00:12:46.40" />
                    <SPLIT distance="1150" swimtime="00:13:21.37" />
                    <SPLIT distance="1200" swimtime="00:13:56.53" />
                    <SPLIT distance="1250" swimtime="00:14:31.15" />
                    <SPLIT distance="1300" swimtime="00:15:06.10" />
                    <SPLIT distance="1350" swimtime="00:15:40.74" />
                    <SPLIT distance="1400" swimtime="00:16:15.29" />
                    <SPLIT distance="1450" swimtime="00:16:50.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1863" points="601" swimtime="00:01:00.31" resultid="5328" heatid="5317" lane="1" entrytime="00:01:00.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:07.11" eventid="1978" heatid="4836" lane="4" />
                <ENTRY entrytime="00:09:09.01" eventid="2020" heatid="4876" lane="4">
                  <MEETINFO qualificationtime="00:09:09.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Tim" gender="M" lastname="Dreher" nation="GER" license="205376" athleteid="3552">
              <RESULTS>
                <RESULT eventid="1749" points="646" swimtime="00:01:54.92" resultid="3553" heatid="4684" lane="4" entrytime="00:01:53.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                    <SPLIT distance="100" swimtime="00:00:56.39" />
                    <SPLIT distance="150" swimtime="00:01:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="543" swimtime="00:02:14.32" resultid="3554" heatid="4755" lane="5" entrytime="00:02:10.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                    <SPLIT distance="100" swimtime="00:01:03.43" />
                    <SPLIT distance="150" swimtime="00:01:44.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:06.68" eventid="2041" heatid="4892" lane="3" />
                <ENTRY entrytime="00:08:53.45" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:08:53.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.92" eventid="1870" heatid="5342" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Luise" gender="F" lastname="Dörries" nation="GER" license="162166" athleteid="3536">
              <RESULTS>
                <RESULT eventid="1771" points="518" swimtime="00:05:22.99" resultid="3537" heatid="4707" lane="3" entrytime="00:05:15.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:10.80" />
                    <SPLIT distance="150" swimtime="00:01:52.33" />
                    <SPLIT distance="200" swimtime="00:02:34.62" />
                    <SPLIT distance="250" swimtime="00:03:22.74" />
                    <SPLIT distance="300" swimtime="00:04:11.71" />
                    <SPLIT distance="350" swimtime="00:04:47.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="647" swimtime="00:04:31.06" resultid="3538" heatid="4763" lane="3" entrytime="00:04:31.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:04.38" />
                    <SPLIT distance="150" swimtime="00:01:38.63" />
                    <SPLIT distance="200" swimtime="00:02:13.06" />
                    <SPLIT distance="250" swimtime="00:02:47.73" />
                    <SPLIT distance="300" swimtime="00:03:22.56" />
                    <SPLIT distance="350" swimtime="00:03:57.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="677" swimtime="00:17:27.04" resultid="3539" heatid="4804" lane="4" entrytime="00:17:32.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="150" swimtime="00:01:42.05" />
                    <SPLIT distance="200" swimtime="00:02:17.36" />
                    <SPLIT distance="250" swimtime="00:02:52.61" />
                    <SPLIT distance="300" swimtime="00:03:27.65" />
                    <SPLIT distance="350" swimtime="00:04:02.87" />
                    <SPLIT distance="400" swimtime="00:04:37.85" />
                    <SPLIT distance="450" swimtime="00:05:12.97" />
                    <SPLIT distance="500" swimtime="00:05:47.83" />
                    <SPLIT distance="550" swimtime="00:06:22.76" />
                    <SPLIT distance="600" swimtime="00:06:57.90" />
                    <SPLIT distance="650" swimtime="00:07:32.78" />
                    <SPLIT distance="700" swimtime="00:08:07.82" />
                    <SPLIT distance="750" swimtime="00:08:42.71" />
                    <SPLIT distance="800" swimtime="00:09:17.74" />
                    <SPLIT distance="850" swimtime="00:09:52.70" />
                    <SPLIT distance="900" swimtime="00:10:27.78" />
                    <SPLIT distance="950" swimtime="00:11:02.81" />
                    <SPLIT distance="1000" swimtime="00:11:37.91" />
                    <SPLIT distance="1050" swimtime="00:12:13.05" />
                    <SPLIT distance="1100" swimtime="00:12:48.04" />
                    <SPLIT distance="1150" swimtime="00:13:23.09" />
                    <SPLIT distance="1200" swimtime="00:13:58.16" />
                    <SPLIT distance="1250" swimtime="00:14:33.28" />
                    <SPLIT distance="1300" swimtime="00:15:08.44" />
                    <SPLIT distance="1350" swimtime="00:15:43.55" />
                    <SPLIT distance="1400" swimtime="00:16:18.53" />
                    <SPLIT distance="1450" swimtime="00:16:53.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.94" eventid="1978" heatid="4838" lane="6" />
                <ENTRY entrytime="00:09:14.39" eventid="2020" heatid="4876" lane="2">
                  <MEETINFO qualificationtime="00:09:14.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Susanne" gender="F" lastname="Dörries" nation="GER" license="157347" athleteid="3542">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.00" eventid="1978" heatid="4836" lane="6" />
                <ENTRY entrytime="NT" eventid="2020" status="RJC" />
                <ENTRY entrytime="00:02:28.00" eventid="2096" heatid="4935" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Dix" gender="M" lastname="Eisenbraun" nation="GER" license="176717" athleteid="3557">
              <RESULTS>
                <RESULT eventid="1763" points="541" swimtime="00:01:08.22" resultid="3558" heatid="4699" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="528" swimtime="00:02:15.60" resultid="3559" heatid="4754" lane="6" entrytime="00:02:14.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="100" swimtime="00:01:04.93" />
                    <SPLIT distance="150" swimtime="00:01:43.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:13.00" eventid="2041" heatid="4892" lane="5" />
                <ENTRY entrytime="00:02:27.00" eventid="2089" heatid="4929" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Sebastian" gender="M" lastname="Greß" nation="GER" license="138833" athleteid="3562">
              <RESULTS>
                <RESULT eventid="1778" points="665" swimtime="00:00:55.47" resultid="3563" heatid="4714" lane="3" entrytime="00:00:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="626" swimtime="00:00:23.68" resultid="3564" heatid="4776" lane="5" entrytime="00:00:24.00" />
                <RESULT eventid="1898" points="672" swimtime="00:00:55.28" resultid="5453" heatid="4717" lane="3" entrytime="00:00:55.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1947" points="624" swimtime="00:00:23.70" resultid="5470" heatid="4778" lane="1" entrytime="00:00:23.68" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:30.00" eventid="1985" heatid="4847" lane="5" />
                <ENTRY entrytime="00:00:59.00" eventid="2027" heatid="4881" lane="4" />
                <ENTRY entrytime="00:00:25.00" eventid="2103" heatid="4947" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lars" gender="M" lastname="Grundheber" nation="GER" license="234237" athleteid="3568">
              <RESULTS>
                <RESULT eventid="1749" points="672" swimtime="00:01:53.41" resultid="3569" heatid="4684" lane="2" entrytime="00:01:53.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.27" />
                    <SPLIT distance="100" swimtime="00:00:54.78" />
                    <SPLIT distance="150" swimtime="00:01:24.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="633" swimtime="00:02:07.67" resultid="3570" heatid="4754" lane="3" entrytime="00:02:05.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="100" swimtime="00:01:01.21" />
                    <SPLIT distance="150" swimtime="00:01:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1926" points="606" swimtime="00:02:09.54" resultid="5434" heatid="4757" lane="1" entrytime="00:02:07.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="100" swimtime="00:01:01.71" />
                    <SPLIT distance="150" swimtime="00:01:39.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:25.52" eventid="1999" heatid="4862" lane="4" />
                <ENTRY entrytime="00:03:59.65" eventid="2075" heatid="4912" lane="5" />
                <ENTRY entrytime="00:08:29.14" eventid="2168" heatid="4809" lane="5">
                  <MEETINFO qualificationtime="00:08:29.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.41" eventid="1870" heatid="4686" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Alina" gender="F" lastname="Hennl" nation="GER" license="173169" athleteid="3574">
              <RESULTS>
                <RESULT eventid="1771" status="DNS" swimtime="00:00:00.00" resultid="3575" heatid="4708" lane="3" entrytime="00:04:54.33" />
                <RESULT eventid="1813" status="DNS" swimtime="00:00:00.00" resultid="3576" heatid="4747" lane="4" entrytime="00:02:18.46" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:09.35" eventid="1978" heatid="4836" lane="2" />
                <ENTRY entrytime="00:02:18.44" eventid="2055" heatid="4902" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Svenja" gender="F" lastname="Herbert" nation="GER" license="304086" athleteid="3579">
              <RESULTS>
                <RESULT eventid="1771" points="591" swimtime="00:05:09.12" resultid="3580" heatid="4708" lane="1" entrytime="00:05:10.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                    <SPLIT distance="150" swimtime="00:01:50.03" />
                    <SPLIT distance="200" swimtime="00:02:29.57" />
                    <SPLIT distance="250" swimtime="00:03:13.21" />
                    <SPLIT distance="300" swimtime="00:03:58.82" />
                    <SPLIT distance="350" swimtime="00:04:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="662" swimtime="00:04:28.99" resultid="3581" heatid="4764" lane="6" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="100" swimtime="00:01:04.40" />
                    <SPLIT distance="150" swimtime="00:01:38.18" />
                    <SPLIT distance="200" swimtime="00:02:12.09" />
                    <SPLIT distance="250" swimtime="00:02:46.44" />
                    <SPLIT distance="300" swimtime="00:03:21.18" />
                    <SPLIT distance="350" swimtime="00:03:55.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="645" swimtime="00:17:44.40" resultid="3582" heatid="4804" lane="1" entrytime="00:17:55.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:05.99" />
                    <SPLIT distance="150" swimtime="00:01:40.67" />
                    <SPLIT distance="200" swimtime="00:02:15.35" />
                    <SPLIT distance="250" swimtime="00:02:50.34" />
                    <SPLIT distance="300" swimtime="00:03:25.52" />
                    <SPLIT distance="350" swimtime="00:04:00.87" />
                    <SPLIT distance="400" swimtime="00:04:36.49" />
                    <SPLIT distance="450" swimtime="00:05:12.30" />
                    <SPLIT distance="500" swimtime="00:05:47.81" />
                    <SPLIT distance="550" swimtime="00:06:23.38" />
                    <SPLIT distance="600" swimtime="00:06:59.11" />
                    <SPLIT distance="650" swimtime="00:07:34.83" />
                    <SPLIT distance="700" swimtime="00:08:10.45" />
                    <SPLIT distance="750" swimtime="00:08:46.25" />
                    <SPLIT distance="800" swimtime="00:09:22.32" />
                    <SPLIT distance="850" swimtime="00:09:58.09" />
                    <SPLIT distance="900" swimtime="00:10:34.07" />
                    <SPLIT distance="950" swimtime="00:11:10.05" />
                    <SPLIT distance="1000" swimtime="00:11:46.09" />
                    <SPLIT distance="1050" swimtime="00:12:21.64" />
                    <SPLIT distance="1100" swimtime="00:12:57.47" />
                    <SPLIT distance="1150" swimtime="00:13:33.75" />
                    <SPLIT distance="1200" swimtime="00:14:09.77" />
                    <SPLIT distance="1250" swimtime="00:14:45.90" />
                    <SPLIT distance="1300" swimtime="00:15:22.07" />
                    <SPLIT distance="1350" swimtime="00:15:57.94" />
                    <SPLIT distance="1400" swimtime="00:16:33.91" />
                    <SPLIT distance="1450" swimtime="00:17:09.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.00" eventid="1978" heatid="4838" lane="5" />
                <ENTRY entrytime="00:02:27.99" eventid="2055" heatid="4902" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Alina" gender="F" lastname="Jungklaus" nation="GER" license="249937" athleteid="3585">
              <RESULTS>
                <RESULT eventid="1059" points="675" swimtime="00:00:58.02" resultid="3586" heatid="4673" lane="3" entrytime="00:00:56.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="748" swimtime="00:04:18.33" resultid="3587" heatid="4764" lane="3" entrytime="00:04:07.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:01:02.16" />
                    <SPLIT distance="150" swimtime="00:01:34.83" />
                    <SPLIT distance="200" swimtime="00:02:07.72" />
                    <SPLIT distance="250" swimtime="00:02:40.76" />
                    <SPLIT distance="300" swimtime="00:03:13.94" />
                    <SPLIT distance="350" swimtime="00:03:47.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="754" swimtime="00:16:50.41" resultid="3588" heatid="4804" lane="3" entrytime="00:16:55.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                    <SPLIT distance="150" swimtime="00:01:37.07" />
                    <SPLIT distance="200" swimtime="00:02:10.72" />
                    <SPLIT distance="250" swimtime="00:02:44.48" />
                    <SPLIT distance="300" swimtime="00:03:18.24" />
                    <SPLIT distance="350" swimtime="00:03:52.20" />
                    <SPLIT distance="400" swimtime="00:04:26.54" />
                    <SPLIT distance="450" swimtime="00:05:00.62" />
                    <SPLIT distance="500" swimtime="00:05:34.57" />
                    <SPLIT distance="550" swimtime="00:06:08.71" />
                    <SPLIT distance="600" swimtime="00:06:42.89" />
                    <SPLIT distance="650" swimtime="00:07:16.92" />
                    <SPLIT distance="700" swimtime="00:07:50.92" />
                    <SPLIT distance="750" swimtime="00:08:24.93" />
                    <SPLIT distance="800" swimtime="00:08:58.86" />
                    <SPLIT distance="850" swimtime="00:09:32.83" />
                    <SPLIT distance="900" swimtime="00:10:06.90" />
                    <SPLIT distance="950" swimtime="00:10:40.91" />
                    <SPLIT distance="1000" swimtime="00:11:15.07" />
                    <SPLIT distance="1050" swimtime="00:11:48.97" />
                    <SPLIT distance="1100" swimtime="00:12:23.09" />
                    <SPLIT distance="1150" swimtime="00:12:57.20" />
                    <SPLIT distance="1200" swimtime="00:13:31.48" />
                    <SPLIT distance="1250" swimtime="00:14:05.01" />
                    <SPLIT distance="1300" swimtime="00:14:39.16" />
                    <SPLIT distance="1350" swimtime="00:15:12.68" />
                    <SPLIT distance="1400" swimtime="00:15:46.51" />
                    <SPLIT distance="1450" swimtime="00:16:19.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:59.16" eventid="1978" heatid="4837" lane="3" />
                <ENTRY entrytime="00:00:27.11" eventid="2082" heatid="4923" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Lena" gender="F" lastname="Kalla" nation="GER" license="143081" athleteid="3591">
              <RESULTS>
                <RESULT eventid="1799" points="628" swimtime="00:01:06.17" resultid="3592" heatid="4734" lane="4" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="648" swimtime="00:00:28.16" resultid="3593" heatid="4800" lane="4" entrytime="00:00:29.00" />
                <RESULT eventid="1919" points="695" swimtime="00:01:03.96" resultid="5392" heatid="4737" lane="3" entrytime="00:01:06.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="631" swimtime="00:00:28.42" resultid="5506" heatid="4802" lane="4" entrytime="00:00:28.16" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.00" eventid="2034" heatid="4888" lane="2" />
                <ENTRY entrytime="00:02:20.00" eventid="2096" heatid="4937" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Jakob" gender="M" lastname="Markowski" nation="GER" license="154737" athleteid="3596">
              <RESULTS>
                <RESULT eventid="1763" points="708" swimtime="00:01:02.39" resultid="3597" heatid="4703" lane="4" entrytime="00:01:03.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="733" swimtime="00:00:22.47" resultid="3598" heatid="4777" lane="3" entrytime="00:00:22.86" />
                <RESULT eventid="1884" points="710" swimtime="00:01:02.31" resultid="5356" heatid="4704" lane="3" entrytime="00:01:02.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1947" points="737" swimtime="00:00:22.42" resultid="5467" heatid="4778" lane="4" entrytime="00:00:22.47" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:28.79" eventid="1985" heatid="4846" lane="3" />
                <ENTRY entrytime="00:00:57.45" eventid="2027" heatid="4881" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Sören" gender="M" lastname="Meißner" nation="GER" license="106221" athleteid="3601">
              <ENTRIES>
                <ENTRY entrytime="00:07:58.29" eventid="2168" heatid="4809" lane="4">
                  <MEETINFO qualificationtime="00:07:58.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Laura" gender="F" lastname="Neumann" nation="GER" license="249654" athleteid="3603">
              <RESULTS>
                <RESULT eventid="1771" points="646" swimtime="00:05:00.13" resultid="3604" heatid="4708" lane="2" entrytime="00:05:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:01:47.42" />
                    <SPLIT distance="200" swimtime="00:02:25.96" />
                    <SPLIT distance="250" swimtime="00:03:08.23" />
                    <SPLIT distance="300" swimtime="00:03:51.27" />
                    <SPLIT distance="350" swimtime="00:04:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1841" points="562" swimtime="00:02:43.04" resultid="3605" heatid="4783" lane="2" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:02:01.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1954" points="566" swimtime="00:02:42.67" resultid="5486" heatid="5491" lane="4" entrytime="00:02:43.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:02:00.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.00" eventid="1978" heatid="4837" lane="5" />
                <ENTRY entrytime="00:02:26.00" eventid="2055" heatid="4903" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Leonie" gender="F" lastname="Neumann" nation="GER" license="249655" athleteid="3608">
              <RESULTS>
                <RESULT eventid="1059" points="579" swimtime="00:01:01.08" resultid="3609" heatid="4674" lane="6" entrytime="00:01:00.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="658" swimtime="00:04:29.58" resultid="3610" heatid="4763" lane="4" entrytime="00:04:32.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                    <SPLIT distance="100" swimtime="00:01:05.14" />
                    <SPLIT distance="150" swimtime="00:01:39.39" />
                    <SPLIT distance="200" swimtime="00:02:13.60" />
                    <SPLIT distance="250" swimtime="00:02:48.20" />
                    <SPLIT distance="300" swimtime="00:03:22.77" />
                    <SPLIT distance="350" swimtime="00:03:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1905" points="652" swimtime="00:17:40.57" resultid="3611" heatid="4804" lane="5" entrytime="00:17:55.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="150" swimtime="00:01:42.38" />
                    <SPLIT distance="200" swimtime="00:02:17.87" />
                    <SPLIT distance="250" swimtime="00:02:53.01" />
                    <SPLIT distance="300" swimtime="00:03:28.30" />
                    <SPLIT distance="350" swimtime="00:04:03.54" />
                    <SPLIT distance="400" swimtime="00:04:38.93" />
                    <SPLIT distance="450" swimtime="00:05:14.37" />
                    <SPLIT distance="500" swimtime="00:05:49.88" />
                    <SPLIT distance="550" swimtime="00:06:25.44" />
                    <SPLIT distance="600" swimtime="00:07:01.26" />
                    <SPLIT distance="650" swimtime="00:07:36.83" />
                    <SPLIT distance="700" swimtime="00:08:12.54" />
                    <SPLIT distance="750" swimtime="00:08:48.24" />
                    <SPLIT distance="800" swimtime="00:09:23.76" />
                    <SPLIT distance="850" swimtime="00:09:59.62" />
                    <SPLIT distance="900" swimtime="00:10:35.22" />
                    <SPLIT distance="950" swimtime="00:11:10.92" />
                    <SPLIT distance="1000" swimtime="00:11:46.43" />
                    <SPLIT distance="1050" swimtime="00:12:21.98" />
                    <SPLIT distance="1100" swimtime="00:12:57.52" />
                    <SPLIT distance="1150" swimtime="00:13:33.13" />
                    <SPLIT distance="1200" swimtime="00:14:08.90" />
                    <SPLIT distance="1250" swimtime="00:14:44.41" />
                    <SPLIT distance="1300" swimtime="00:15:20.15" />
                    <SPLIT distance="1350" swimtime="00:15:55.51" />
                    <SPLIT distance="1400" swimtime="00:16:30.94" />
                    <SPLIT distance="1450" swimtime="00:17:05.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:10.00" eventid="1978" heatid="4836" lane="5" />
                <ENTRY entrytime="00:09:23.26" eventid="2020" heatid="4876" lane="1">
                  <MEETINFO qualificationtime="00:09:19.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Natalie" gender="F" lastname="Schnabel" nation="GER" license="299453" athleteid="3614">
              <RESULTS>
                <RESULT eventid="1059" points="539" swimtime="00:01:02.52" resultid="3615" heatid="4665" lane="1" entrytime="00:01:03.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="494" swimtime="00:00:36.43" resultid="3616" heatid="4688" lane="1" entrytime="00:00:37.43" />
                <RESULT eventid="1841" points="480" swimtime="00:02:51.82" resultid="3617" heatid="4780" lane="6" entrytime="00:02:55.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:06.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:18.78" eventid="1992" heatid="4853" lane="2" />
                <ENTRY entrytime="00:02:35.06" eventid="2055" heatid="4900" lane="5" />
                <ENTRY entrytime="00:00:29.00" eventid="2082" heatid="4917" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Ruwen" gender="M" lastname="Straub" nation="GER" license="148906" athleteid="3621">
              <RESULTS>
                <RESULT eventid="1749" points="686" swimtime="00:01:52.64" resultid="3622" heatid="4685" lane="4" entrytime="00:01:51.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                    <SPLIT distance="100" swimtime="00:00:55.22" />
                    <SPLIT distance="150" swimtime="00:01:23.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="531" swimtime="00:02:10.44" resultid="3623" heatid="4789" lane="6" entrytime="00:02:17.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="100" swimtime="00:01:03.81" />
                    <SPLIT distance="150" swimtime="00:01:37.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:52.90" eventid="1971" heatid="4827" lane="5" />
                <ENTRY entrytime="00:03:45.56" eventid="2075" heatid="4912" lane="3" />
                <ENTRY entrytime="00:07:54.96" eventid="2168" heatid="4809" lane="3">
                  <MEETINFO qualificationtime="00:07:54.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.64" eventid="1870" heatid="4686" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Shay" gender="M" lastname="Toledano" nation="GER" license="365525" athleteid="3627">
              <RESULTS>
                <RESULT eventid="1792" points="692" swimtime="00:15:58.60" resultid="3628" heatid="4727" lane="3" entrytime="00:15:48.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:33.00" />
                    <SPLIT distance="200" swimtime="00:02:04.42" />
                    <SPLIT distance="250" swimtime="00:02:35.81" />
                    <SPLIT distance="300" swimtime="00:03:07.47" />
                    <SPLIT distance="350" swimtime="00:03:39.12" />
                    <SPLIT distance="400" swimtime="00:04:10.78" />
                    <SPLIT distance="450" swimtime="00:04:42.61" />
                    <SPLIT distance="500" swimtime="00:05:14.43" />
                    <SPLIT distance="550" swimtime="00:05:46.46" />
                    <SPLIT distance="600" swimtime="00:06:18.76" />
                    <SPLIT distance="650" swimtime="00:06:50.44" />
                    <SPLIT distance="700" swimtime="00:07:22.52" />
                    <SPLIT distance="750" swimtime="00:07:54.59" />
                    <SPLIT distance="800" swimtime="00:08:26.66" />
                    <SPLIT distance="850" swimtime="00:08:58.79" />
                    <SPLIT distance="900" swimtime="00:09:31.19" />
                    <SPLIT distance="950" swimtime="00:10:03.22" />
                    <SPLIT distance="1000" swimtime="00:10:35.46" />
                    <SPLIT distance="1050" swimtime="00:11:07.94" />
                    <SPLIT distance="1100" swimtime="00:11:40.34" />
                    <SPLIT distance="1150" swimtime="00:12:12.83" />
                    <SPLIT distance="1200" swimtime="00:12:45.10" />
                    <SPLIT distance="1250" swimtime="00:13:17.32" />
                    <SPLIT distance="1300" swimtime="00:13:49.55" />
                    <SPLIT distance="1350" swimtime="00:14:21.87" />
                    <SPLIT distance="1400" swimtime="00:14:54.51" />
                    <SPLIT distance="1450" swimtime="00:15:27.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:45.03" eventid="1999" heatid="4861" lane="3" />
                <ENTRY entrytime="00:04:08.47" eventid="2075" heatid="4911" lane="2" />
                <ENTRY entrytime="00:08:47.66" eventid="2168" heatid="4808" lane="1">
                  <MEETINFO qualificationtime="00:08:47.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Svenja" gender="F" lastname="Zihsler" nation="GER" license="151222" athleteid="3632">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.52" eventid="1978" heatid="4836" lane="3" />
                <ENTRY entrytime="00:08:40.16" eventid="2020" heatid="4876" lane="3">
                  <MEETINFO qualificationtime="00:08:40.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.74" eventid="2055" heatid="4903" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="2048" points="679" swimtime="00:01:42.97" resultid="3636" heatid="4806" lane="4" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                    <SPLIT distance="100" swimtime="00:00:56.23" />
                    <SPLIT distance="150" swimtime="00:01:21.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3497" number="1" />
                    <RELAYPOSITION athleteid="3524" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="3562" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="3596" number="4" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:26.89" eventid="2232" heatid="4812" lane="3" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="2062" points="701" swimtime="00:01:57.08" resultid="3638" heatid="4807" lane="4" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                    <SPLIT distance="100" swimtime="00:01:01.95" />
                    <SPLIT distance="150" swimtime="00:01:30.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3591" number="1" />
                    <RELAYPOSITION athleteid="3502" number="2" />
                    <RELAYPOSITION athleteid="3530" number="3" />
                    <RELAYPOSITION athleteid="3585" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:47.00" eventid="2224" heatid="4810" lane="4" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5806" nation="GER" region="02" clubid="2708" name="Team Buron Kaufbeuren">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Nadja" gender="F" lastname="Amrhein" nation="GER" license="262168" swrid="4491234" athleteid="2709">
              <ENTRIES>
                <ENTRY entrytime="00:01:17.55" eventid="1992" heatid="4854" lane="6" />
                <ENTRY entrytime="00:02:32.52" eventid="2055" heatid="4902" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Katharina" gender="F" lastname="Breunig" nation="GER" license="299621" athleteid="2712">
              <RESULTS>
                <RESULT eventid="1059" points="472" swimtime="00:01:05.37" resultid="2713" heatid="4663" lane="5" entrytime="00:01:04.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1756" points="420" swimtime="00:00:38.43" resultid="2714" heatid="4687" lane="4" entrytime="00:00:37.66" />
                <RESULT eventid="1785" points="428" swimtime="00:01:12.97" resultid="2715" heatid="4719" lane="2" entrytime="00:01:12.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="459" swimtime="00:01:13.43" resultid="2716" heatid="4732" lane="3" entrytime="00:01:12.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:20.16" eventid="1978" heatid="4830" lane="2" />
                <ENTRY entrytime="00:00:33.91" eventid="2034" heatid="4884" lane="2" />
                <ENTRY entrytime="00:02:38.37" eventid="2055" heatid="4898" lane="1" />
                <ENTRY entrytime="00:02:33.79" eventid="2096" heatid="4933" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Gina" gender="F" lastname="Mayer" nation="GER" license="257249" athleteid="2721">
              <RESULTS>
                <RESULT eventid="1059" points="522" swimtime="00:01:03.21" resultid="2722" heatid="4670" lane="6" entrytime="00:01:02.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="450" swimtime="00:01:13.92" resultid="2723" heatid="4733" lane="4" entrytime="00:01:11.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="500" swimtime="00:04:55.35" resultid="2724" heatid="4761" lane="6" entrytime="00:04:48.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:44.40" />
                    <SPLIT distance="200" swimtime="00:02:21.87" />
                    <SPLIT distance="250" swimtime="00:03:00.11" />
                    <SPLIT distance="300" swimtime="00:03:38.59" />
                    <SPLIT distance="350" swimtime="00:04:17.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:12.97" eventid="1978" heatid="4835" lane="1" />
                <ENTRY entrytime="00:00:32.66" eventid="2034" heatid="4886" lane="2" />
                <ENTRY entrytime="00:02:34.12" eventid="2055" heatid="4901" lane="6" />
                <ENTRY entrytime="00:00:28.84" eventid="2082" heatid="4918" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Wolfgang" gender="M" lastname="Orth" nation="GER" license="226633" athleteid="2729">
              <RESULTS>
                <RESULT eventid="1749" points="562" swimtime="00:02:00.35" resultid="2730" heatid="4683" lane="6" entrytime="00:01:58.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                    <SPLIT distance="100" swimtime="00:00:58.48" />
                    <SPLIT distance="150" swimtime="00:01:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1792" points="595" swimtime="00:16:48.21" resultid="2731" heatid="4727" lane="2" entrytime="00:16:27.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                    <SPLIT distance="100" swimtime="00:01:01.92" />
                    <SPLIT distance="150" swimtime="00:01:35.27" />
                    <SPLIT distance="200" swimtime="00:02:08.49" />
                    <SPLIT distance="250" swimtime="00:02:41.91" />
                    <SPLIT distance="300" swimtime="00:03:15.25" />
                    <SPLIT distance="350" swimtime="00:03:48.75" />
                    <SPLIT distance="400" swimtime="00:04:22.62" />
                    <SPLIT distance="450" swimtime="00:04:56.44" />
                    <SPLIT distance="500" swimtime="00:05:30.26" />
                    <SPLIT distance="550" swimtime="00:06:03.96" />
                    <SPLIT distance="600" swimtime="00:06:37.80" />
                    <SPLIT distance="650" swimtime="00:07:11.96" />
                    <SPLIT distance="700" swimtime="00:07:45.82" />
                    <SPLIT distance="750" swimtime="00:08:19.58" />
                    <SPLIT distance="800" swimtime="00:08:53.79" />
                    <SPLIT distance="850" swimtime="00:09:28.32" />
                    <SPLIT distance="900" swimtime="00:10:02.29" />
                    <SPLIT distance="950" swimtime="00:10:36.25" />
                    <SPLIT distance="1000" swimtime="00:11:10.20" />
                    <SPLIT distance="1050" swimtime="00:11:44.20" />
                    <SPLIT distance="1100" swimtime="00:12:18.29" />
                    <SPLIT distance="1150" swimtime="00:12:52.05" />
                    <SPLIT distance="1200" swimtime="00:13:26.16" />
                    <SPLIT distance="1250" swimtime="00:14:00.14" />
                    <SPLIT distance="1300" swimtime="00:14:34.05" />
                    <SPLIT distance="1350" swimtime="00:15:08.00" />
                    <SPLIT distance="1400" swimtime="00:15:42.04" />
                    <SPLIT distance="1450" swimtime="00:16:15.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="425" swimtime="00:02:20.43" resultid="2732" heatid="4790" lane="6" entrytime="00:02:15.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:44.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:55.62" eventid="1971" heatid="4821" lane="5" />
                <ENTRY entrytime="00:01:03.56" eventid="2013" heatid="4870" lane="2" />
                <ENTRY entrytime="00:04:11.03" eventid="2075" heatid="4911" lane="6" />
                <ENTRY entrytime="00:08:48.98" eventid="2168" heatid="4808" lane="6">
                  <MEETINFO qualificationtime="00:08:48.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Johannes" gender="M" lastname="Vorbach" nation="GER" license="257156" athleteid="2737">
              <RESULTS>
                <RESULT eventid="1763" points="428" swimtime="00:01:13.76" resultid="2738" heatid="4696" lane="3" entrytime="00:01:13.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="419" swimtime="00:00:27.07" resultid="2739" heatid="4765" lane="4" entrytime="00:00:27.37" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.81" eventid="1971" heatid="4815" lane="6" />
                <ENTRY entrytime="00:00:33.61" eventid="1985" heatid="4842" lane="6" />
                <ENTRY entrytime="00:02:42.43" eventid="2089" heatid="4925" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Lea" gender="F" lastname="Wienstruck" nation="GER" license="296635" athleteid="2743">
              <RESULTS>
                <RESULT eventid="1059" points="517" swimtime="00:01:03.41" resultid="2744" heatid="4664" lane="4" entrytime="00:01:03.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="470" swimtime="00:01:10.77" resultid="2745" heatid="4721" lane="1" entrytime="00:01:10.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="493" swimtime="00:01:11.71" resultid="2746" heatid="4733" lane="1" entrytime="00:01:12.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.59" eventid="2034" heatid="4886" lane="4" />
                <ENTRY entrytime="00:02:34.66" eventid="2055" heatid="4900" lane="3" />
                <ENTRY entrytime="00:00:29.22" eventid="2082" heatid="4916" lane="5" />
                <ENTRY entrytime="00:02:29.99" eventid="2096" heatid="4934" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4397" nation="GER" region="02" clubid="2751" name="TG Kitzingen">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Viktoria" gender="F" lastname="Kolb" nation="GER" license="291280" athleteid="2752">
              <RESULTS>
                <RESULT eventid="1059" points="488" swimtime="00:01:04.66" resultid="2753" heatid="4665" lane="3" entrytime="00:01:03.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="421" swimtime="00:01:15.57" resultid="2754" heatid="4729" lane="2" entrytime="00:01:14.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4405" nation="GER" region="02" clubid="4159" name="TSG Kleinostheim">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Francis" gender="M" lastname="Hartl" nation="GER" license="285486" athleteid="4163">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.09" eventid="1971" heatid="4813" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Alena" gender="F" lastname="Hennl" nation="GER" license="208754" athleteid="4165">
              <RESULTS>
                <RESULT eventid="1756" points="630" swimtime="00:00:33.58" resultid="4166" heatid="4693" lane="2" entrytime="00:00:33.93" />
                <RESULT eventid="1813" points="514" swimtime="00:02:29.26" resultid="4167" heatid="4747" lane="2" entrytime="00:02:25.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:09.82" />
                    <SPLIT distance="150" swimtime="00:01:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="560" swimtime="00:00:29.57" resultid="4168" heatid="4801" lane="6" entrytime="00:00:29.91" />
                <RESULT eventid="1877" points="638" swimtime="00:00:33.44" resultid="5346" heatid="4695" lane="5" entrytime="00:00:33.58" />
                <RESULT eventid="1933" points="505" swimtime="00:02:30.11" resultid="5424" heatid="5429" lane="3" entrytime="00:02:29.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:50.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="547" swimtime="00:00:29.80" resultid="5512" heatid="5517" lane="4" entrytime="00:00:29.57" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:16.85" eventid="1992" heatid="4855" lane="6" />
                <ENTRY entrytime="00:01:05.46" eventid="2006" heatid="4866" lane="2" />
                <ENTRY entrytime="00:02:28.56" eventid="2055" heatid="4902" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4439" nation="GER" region="02" clubid="2481" name="TSV - Eintracht Karlsfeld">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Johannes" gender="M" lastname="Heizenreder" nation="GER" license="248442" athleteid="2482">
              <RESULTS>
                <RESULT eventid="1806" points="378" swimtime="00:00:30.73" resultid="2483" heatid="4741" lane="6" entrytime="00:00:29.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Miriam" gender="F" lastname="Zanklmaier" nation="GER" license="283818" athleteid="2484">
              <RESULTS>
                <RESULT eventid="1756" points="500" swimtime="00:00:36.27" resultid="2485" heatid="4690" lane="6" entrytime="00:00:36.50" />
                <RESULT eventid="1799" points="501" swimtime="00:01:11.31" resultid="2486" heatid="4734" lane="1" entrytime="00:01:11.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="512" swimtime="00:00:30.47" resultid="2487" heatid="4799" lane="2" entrytime="00:00:30.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4413" nation="GER" region="02" clubid="2674" name="TSV 1860 Rosenheim">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Alexander" gender="M" lastname="Bauer" nation="GER" license="257560" athleteid="2675">
              <RESULTS>
                <RESULT eventid="1778" points="455" swimtime="00:01:02.97" resultid="2676" heatid="4711" lane="6" entrytime="00:01:02.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:28.45" eventid="2103" heatid="4941" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Paula" gender="F" lastname="Borst" nation="GER" license="200640" athleteid="2678">
              <RESULTS>
                <RESULT eventid="1059" points="527" swimtime="00:01:03.00" resultid="2679" heatid="4670" lane="5" entrytime="00:01:01.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="474" swimtime="00:00:31.25" resultid="2680" heatid="4799" lane="4" entrytime="00:00:30.50" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:28.20" eventid="2082" heatid="4922" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lucas" gender="M" lastname="Kleinicke" nation="GER" license="226836" athleteid="2682">
              <RESULTS>
                <RESULT eventid="1749" points="438" swimtime="00:02:10.75" resultid="2683" heatid="4678" lane="1" entrytime="00:02:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                    <SPLIT distance="150" swimtime="00:01:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="475" swimtime="00:01:02.08" resultid="2684" heatid="4712" lane="4" entrytime="00:01:01.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="525" swimtime="00:00:25.11" resultid="2685" heatid="4774" lane="5" entrytime="00:00:24.86" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.20" eventid="1971" heatid="4818" lane="6" />
                <ENTRY entrytime="00:00:27.42" eventid="2103" heatid="4943" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Alexandra" gender="F" lastname="Schöne" nation="GER" license="266174" athleteid="2688">
              <RESULTS>
                <RESULT eventid="1059" points="539" swimtime="00:01:02.52" resultid="2689" heatid="4669" lane="3" entrytime="00:01:02.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="471" swimtime="00:01:10.69" resultid="2690" heatid="4721" lane="3" entrytime="00:01:08.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="542" swimtime="00:04:47.57" resultid="2691" heatid="4762" lane="5" entrytime="00:04:41.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                    <SPLIT distance="150" swimtime="00:01:45.42" />
                    <SPLIT distance="200" swimtime="00:02:22.40" />
                    <SPLIT distance="250" swimtime="00:02:59.55" />
                    <SPLIT distance="300" swimtime="00:03:36.31" />
                    <SPLIT distance="350" swimtime="00:04:12.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:12.25" eventid="1978" heatid="4835" lane="4" />
                <ENTRY entrytime="00:00:30.90" eventid="2034" heatid="4889" lane="2" />
                <ENTRY entrytime="00:00:28.30" eventid="2082" heatid="4920" lane="2" />
                <ENTRY entrytime="00:02:33.62" eventid="2096" heatid="4933" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Sarah" gender="F" lastname="Wieser" nation="GER" license="295252" athleteid="2696">
              <RESULTS>
                <RESULT eventid="1855" points="440" swimtime="00:00:32.03" resultid="2697" heatid="4794" lane="5" entrytime="00:00:32.07" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:34.27" eventid="2034" heatid="4883" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4441" nation="GER" region="02" clubid="3253" name="TSV Erding">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Carina" gender="F" lastname="Michaelis" nation="GER" license="313153" athleteid="3254">
              <RESULTS>
                <RESULT eventid="1059" points="526" swimtime="00:01:03.04" resultid="3255" heatid="4666" lane="3" entrytime="00:01:03.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="492" swimtime="00:01:11.78" resultid="3256" heatid="4732" lane="6" entrytime="00:01:12.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="529" swimtime="00:04:49.96" resultid="3257" heatid="4758" lane="3" entrytime="00:04:55.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                    <SPLIT distance="150" swimtime="00:01:44.84" />
                    <SPLIT distance="200" swimtime="00:02:21.94" />
                    <SPLIT distance="250" swimtime="00:02:59.15" />
                    <SPLIT distance="300" swimtime="00:03:36.53" />
                    <SPLIT distance="350" swimtime="00:04:13.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="519" swimtime="00:00:30.33" resultid="3258" heatid="4799" lane="1" entrytime="00:00:30.67" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:15.65" eventid="1978" heatid="4833" lane="5" />
                <ENTRY entrytime="00:00:33.97" eventid="2034" heatid="4884" lane="5" />
                <ENTRY entrytime="00:02:37.06" eventid="2055" heatid="4899" lane="1" />
                <ENTRY entrytime="00:00:28.97" eventid="2082" heatid="4917" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4452" nation="GER" region="02" clubid="2771" name="TSV Hohenbrunn-Riemerl.">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Nick" gender="M" lastname="Bongartz" nation="GER" license="325785" athleteid="2772">
              <RESULTS>
                <RESULT eventid="1749" points="525" swimtime="00:02:03.15" resultid="2773" heatid="4679" lane="5" entrytime="00:02:05.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="100" swimtime="00:01:00.10" />
                    <SPLIT distance="150" swimtime="00:01:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="500" swimtime="00:02:18.11" resultid="2774" heatid="4752" lane="1" entrytime="00:02:20.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:46.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.45" eventid="1971" heatid="4817" lane="4" />
                <ENTRY entrytime="00:05:02.54" eventid="1999" heatid="4860" lane="2" />
                <ENTRY entrytime="00:04:33.74" eventid="2075" heatid="4908" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Adrien" gender="M" lastname="Cara" nation="GER" license="294598" athleteid="2778">
              <RESULTS>
                <RESULT eventid="1763" points="450" swimtime="00:01:12.56" resultid="2779" heatid="4697" lane="5" entrytime="00:01:13.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="496" swimtime="00:02:18.45" resultid="2780" heatid="4750" lane="3" entrytime="00:02:22.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:04.90" />
                    <SPLIT distance="150" swimtime="00:01:45.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="459" swimtime="00:02:16.91" resultid="2781" heatid="4788" lane="3" entrytime="00:02:17.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:05.97" />
                    <SPLIT distance="150" swimtime="00:01:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="460" swimtime="00:02:16.77" resultid="5503" heatid="5504" lane="6" entrytime="00:02:16.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.20" />
                    <SPLIT distance="100" swimtime="00:01:06.13" />
                    <SPLIT distance="150" swimtime="00:01:42.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.50" eventid="1971" heatid="4817" lane="2" />
                <ENTRY entrytime="00:04:59.19" eventid="1999" heatid="4860" lane="4" />
                <ENTRY entrytime="00:01:03.36" eventid="2013" heatid="4870" lane="3" />
                <ENTRY entrytime="00:02:38.40" eventid="2089" heatid="4926" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Daniela" gender="F" lastname="Ernst" nation="GER" license="316890" athleteid="2786">
              <RESULTS>
                <RESULT eventid="1785" points="501" swimtime="00:01:09.25" resultid="2787" heatid="4720" lane="1" entrytime="00:01:11.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:33.98" eventid="2034" heatid="4884" lane="1" />
                <ENTRY entrytime="00:02:32.23" eventid="2096" heatid="4934" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lisa-Marie" gender="F" lastname="Geisler" nation="GER" license="221272" athleteid="2790">
              <RESULTS>
                <RESULT eventid="1756" points="483" swimtime="00:00:36.70" resultid="2791" heatid="4690" lane="4" entrytime="00:00:36.03" />
                <RESULT eventid="1841" points="486" swimtime="00:02:51.14" resultid="2792" heatid="4781" lane="4" entrytime="00:02:49.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:22.55" />
                    <SPLIT distance="150" swimtime="00:02:07.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:17.28" eventid="1992" heatid="4854" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Amna" gender="F" lastname="Hasanbegovic" nation="GER" license="225371" athleteid="2794">
              <RESULTS>
                <RESULT eventid="1799" points="475" swimtime="00:01:12.59" resultid="2795" heatid="4731" lane="4" entrytime="00:01:12.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="497" swimtime="00:00:30.76" resultid="2796" heatid="4797" lane="1" entrytime="00:00:31.08" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:08.34" eventid="2006" heatid="4865" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Eric Florian" gender="M" lastname="Henschel" nation="GER" license="212691" athleteid="2798">
              <RESULTS>
                <RESULT eventid="1834" points="584" swimtime="00:00:24.23" resultid="2799" heatid="4771" lane="1" entrytime="00:00:25.66" />
                <RESULT eventid="1947" points="588" swimtime="00:00:24.18" resultid="5476" heatid="5478" lane="1" entrytime="00:00:24.23" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.98" eventid="1971" heatid="4818" lane="5" />
                <ENTRY entrytime="00:00:27.42" eventid="2103" heatid="4943" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Alina" gender="F" lastname="Hermeking" nation="GER" license="290265" athleteid="2802">
              <RESULTS>
                <RESULT eventid="1756" points="471" swimtime="00:00:36.99" resultid="2803" heatid="4688" lane="2" entrytime="00:00:37.33" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:22.48" eventid="1992" heatid="4850" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Fabian" gender="M" lastname="Hoffmann" nation="GER" license="290269" athleteid="2805">
              <RESULTS>
                <RESULT eventid="1806" points="402" swimtime="00:00:30.10" resultid="2806" heatid="4738" lane="3" entrytime="00:00:31.05" />
                <RESULT eventid="1834" points="440" swimtime="00:00:26.62" resultid="2807" heatid="4768" lane="1" entrytime="00:00:26.46" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:59.46" eventid="1971" heatid="4814" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Tobias" gender="M" lastname="Hollaus" nation="GER" license="209181" athleteid="2809">
              <RESULTS>
                <RESULT eventid="1763" points="652" swimtime="00:01:04.10" resultid="2810" heatid="4702" lane="2" entrytime="00:01:04.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1884" points="676" swimtime="00:01:03.34" resultid="5360" heatid="4704" lane="1" entrytime="00:01:04.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.90" eventid="1985" heatid="4848" lane="5" />
                <ENTRY entrytime="00:02:22.45" eventid="2089" heatid="4928" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Sarah-Isabelle" gender="F" lastname="Mai" nation="GER" license="269795" athleteid="2813">
              <RESULTS>
                <RESULT eventid="1756" points="563" swimtime="00:00:34.86" resultid="2814" heatid="4693" lane="5" entrytime="00:00:34.56" />
                <RESULT eventid="1799" points="503" swimtime="00:01:11.25" resultid="2815" heatid="4736" lane="5" entrytime="00:01:09.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="(Zeit: 14:42), Die Schwimmerin hat bei der 175m Wende nicht mit beiden Händen gleichzeitig angeschlagen" eventid="1841" status="DSQ" swimtime="00:02:47.89" resultid="2816" heatid="4783" lane="1" entrytime="00:02:45.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                    <SPLIT distance="150" swimtime="00:02:03.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:15.81" eventid="1992" heatid="4856" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Francesco" gender="M" lastname="Montanari" nation="GER" license="281775" athleteid="2818">
              <RESULTS>
                <RESULT eventid="1834" points="551" swimtime="00:00:24.71" resultid="2819" heatid="4773" lane="3" entrytime="00:00:24.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Tom" gender="M" lastname="Nolte" nation="GER" license="288931" athleteid="2820">
              <RESULTS>
                <RESULT eventid="1763" points="502" swimtime="00:01:09.94" resultid="2821" heatid="4698" lane="6" entrytime="00:01:11.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="437" swimtime="00:00:29.26" resultid="2822" heatid="4739" lane="3" entrytime="00:00:30.16" />
                <RESULT eventid="1834" points="474" swimtime="00:00:25.97" resultid="2823" heatid="4770" lane="2" entrytime="00:00:25.92" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.81" eventid="1985" heatid="4842" lane="2" />
                <ENTRY entrytime="00:01:06.15" eventid="2013" heatid="4869" lane="2" />
                <ENTRY entrytime="00:00:28.85" eventid="2103" heatid="4940" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Sven" gender="M" lastname="Pesut" nation="GER" license="360757" athleteid="2827">
              <RESULTS>
                <RESULT eventid="1749" points="526" swimtime="00:02:03.07" resultid="2828" heatid="4680" lane="6" entrytime="00:02:04.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="100" swimtime="00:00:59.41" />
                    <SPLIT distance="150" swimtime="00:01:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="488" swimtime="00:01:01.50" resultid="2829" heatid="4712" lane="6" entrytime="00:01:01.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="493" swimtime="00:02:18.75" resultid="2830" heatid="4751" lane="1" entrytime="00:02:22.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                    <SPLIT distance="150" swimtime="00:01:45.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.72" eventid="1971" heatid="4819" lane="3" />
                <ENTRY entrytime="00:05:06.39" eventid="1999" heatid="4859" lane="4" />
                <ENTRY entrytime="00:04:31.63" eventid="2075" heatid="4908" lane="2" />
                <ENTRY entrytime="00:00:27.56" eventid="2103" heatid="4943" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Noah" gender="M" lastname="Rueff" nation="GER" license="241485" athleteid="2835">
              <RESULTS>
                <RESULT eventid="1778" points="444" swimtime="00:01:03.47" resultid="2836" heatid="4710" lane="3" entrytime="00:01:02.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="403" swimtime="00:00:30.07" resultid="2837" heatid="4739" lane="2" entrytime="00:00:30.30" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:33.00" eventid="1985" heatid="4842" lane="5" />
                <ENTRY entrytime="00:01:05.20" eventid="2013" heatid="4869" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Moritz" gender="M" lastname="Schepp" nation="GER" license="279390" athleteid="2840">
              <RESULTS>
                <RESULT eventid="1806" points="437" swimtime="00:00:29.28" resultid="2841" heatid="4739" lane="4" entrytime="00:00:30.27" />
                <RESULT eventid="1834" points="488" swimtime="00:00:25.72" resultid="2842" heatid="4768" lane="2" entrytime="00:00:26.33" />
                <RESULT eventid="1848" points="447" swimtime="00:02:18.14" resultid="2843" heatid="4787" lane="4" entrytime="00:02:20.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:42.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.07" eventid="1971" heatid="4816" lane="1" />
                <ENTRY entrytime="00:01:06.39" eventid="2013" heatid="4869" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Florian" gender="M" lastname="Schimanski" nation="GER" license="183469" athleteid="2846">
              <RESULTS>
                <RESULT eventid="1778" points="523" swimtime="00:01:00.12" resultid="2847" heatid="4713" lane="4" entrytime="00:01:00.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="507" swimtime="00:00:25.40" resultid="2848" heatid="4774" lane="6" entrytime="00:00:24.94" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.07" eventid="1971" heatid="4824" lane="2" />
                <ENTRY entrytime="00:00:25.60" eventid="2103" heatid="4947" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Nico" gender="M" lastname="Schmid" nation="GER" license="175732" athleteid="2851">
              <RESULTS>
                <RESULT eventid="1749" points="608" swimtime="00:01:57.24" resultid="2852" heatid="4685" lane="6" entrytime="00:01:57.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                    <SPLIT distance="100" swimtime="00:00:56.57" />
                    <SPLIT distance="150" swimtime="00:01:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="582" swimtime="00:02:11.29" resultid="2853" heatid="4755" lane="2" entrytime="00:02:09.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="100" swimtime="00:01:02.82" />
                    <SPLIT distance="150" swimtime="00:01:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="553" swimtime="00:00:24.67" resultid="2854" heatid="4775" lane="6" entrytime="00:00:24.63" />
                <RESULT eventid="1926" points="587" swimtime="00:02:10.93" resultid="5440" heatid="5442" lane="1" entrytime="00:02:11.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="100" swimtime="00:01:03.23" />
                    <SPLIT distance="150" swimtime="00:01:41.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:04:35.89" eventid="1999" heatid="4862" lane="2" />
                <ENTRY entrytime="00:04:08.23" eventid="2075" heatid="4911" lane="4" />
                <ENTRY entrytime="NT" eventid="2168" status="RJC" />
                <ENTRY entrytime="00:01:57.24" eventid="1870" heatid="5342" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Magnus" gender="M" lastname="Schweiger" nation="GER" license="158545" athleteid="2858">
              <RESULTS>
                <RESULT eventid="1749" points="661" swimtime="00:01:54.03" resultid="2859" heatid="4685" lane="2" entrytime="00:01:53.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="100" swimtime="00:00:55.26" />
                    <SPLIT distance="150" swimtime="00:01:24.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="584" swimtime="00:00:57.93" resultid="2860" heatid="4716" lane="5" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1898" points="548" swimtime="00:00:59.16" resultid="5456" heatid="4717" lane="5" entrytime="00:00:57.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:53.55" eventid="1971" heatid="4826" lane="6" />
                <ENTRY entrytime="00:02:10.69" eventid="2041" heatid="4893" lane="2" />
                <ENTRY entrytime="00:04:03.77" eventid="2075" heatid="4912" lane="6" />
                <ENTRY entrytime="00:01:54.03" eventid="1870" heatid="4686" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Helena" gender="F" lastname="Sedlar" nation="GER" license="290267" athleteid="2864">
              <RESULTS>
                <RESULT eventid="1059" points="510" swimtime="00:01:03.68" resultid="2865" heatid="4667" lane="5" entrytime="00:01:02.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="532" swimtime="00:04:49.38" resultid="2866" heatid="4759" lane="1" entrytime="00:04:55.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:47.21" />
                    <SPLIT distance="200" swimtime="00:02:24.36" />
                    <SPLIT distance="250" swimtime="00:03:01.44" />
                    <SPLIT distance="300" swimtime="00:03:38.29" />
                    <SPLIT distance="350" swimtime="00:04:15.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="429" swimtime="00:00:32.32" resultid="2867" heatid="4795" lane="1" entrytime="00:00:31.78" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:21.10" eventid="1978" heatid="4829" lane="2" />
                <ENTRY entrytime="00:00:30.03" eventid="2082" heatid="4913" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lana" gender="F" lastname="Sokac" nation="GER" license="360313" athleteid="2870">
              <RESULTS>
                <RESULT eventid="1059" points="643" swimtime="00:00:58.97" resultid="2871" heatid="4674" lane="2" entrytime="00:00:58.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="593" swimtime="00:01:07.42" resultid="2872" heatid="4736" lane="2" entrytime="00:01:07.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="599" swimtime="00:00:28.92" resultid="2873" heatid="4801" lane="2" entrytime="00:00:29.35" />
                <RESULT eventid="1863" points="666" swimtime="00:00:58.29" resultid="5319" heatid="4675" lane="4" entrytime="00:00:58.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1919" points="597" swimtime="00:01:07.27" resultid="5396" heatid="4737" lane="1" entrytime="00:01:07.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1940" points="599" swimtime="00:00:28.91" resultid="5508" heatid="4802" lane="5" entrytime="00:00:28.92" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:06.20" eventid="2006" heatid="4867" lane="5" />
                <ENTRY entrytime="00:00:26.68" eventid="2082" heatid="4922" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Jacopo" gender="M" lastname="Vercelli" nation="GER" license="329282" athleteid="2876">
              <RESULTS>
                <RESULT eventid="1778" points="450" swimtime="00:01:03.18" resultid="2877" heatid="4709" lane="5" entrytime="00:01:04.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="441" swimtime="00:00:26.61" resultid="2878" heatid="4767" lane="4" entrytime="00:00:26.70" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.50" eventid="1971" heatid="4815" lane="5" />
                <ENTRY entrytime="00:02:24.00" eventid="2041" heatid="4891" lane="2" />
                <ENTRY entrytime="00:00:29.00" eventid="2103" heatid="4939" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Sina" gender="F" lastname="Wappenschmidt" nation="GER" license="269801" swrid="4642730" athleteid="2882">
              <RESULTS>
                <RESULT eventid="1059" points="539" swimtime="00:01:02.54" resultid="2883" heatid="4667" lane="3" entrytime="00:01:02.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1785" points="488" swimtime="00:01:09.89" resultid="2884" heatid="4720" lane="4" entrytime="00:01:10.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="598" swimtime="00:04:38.36" resultid="2885" heatid="4761" lane="5" entrytime="00:04:46.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:42.58" />
                    <SPLIT distance="200" swimtime="00:02:18.33" />
                    <SPLIT distance="250" swimtime="00:02:53.80" />
                    <SPLIT distance="300" swimtime="00:03:29.29" />
                    <SPLIT distance="350" swimtime="00:04:04.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:17.63" eventid="1978" heatid="4832" lane="1" />
                <ENTRY entrytime="00:02:33.79" eventid="2055" heatid="4901" lane="2" />
                <ENTRY entrytime="00:02:33.74" eventid="2096" heatid="4933" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Florian" gender="M" lastname="Wutz" nation="GER" license="233903" athleteid="2890">
              <RESULTS>
                <RESULT eventid="1749" points="543" swimtime="00:02:01.73" resultid="2891" heatid="4681" lane="2" entrytime="00:02:02.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="100" swimtime="00:00:59.31" />
                    <SPLIT distance="150" swimtime="00:01:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="530" swimtime="00:00:25.02" resultid="2892" heatid="4769" lane="5" entrytime="00:00:26.17" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.34" eventid="1971" heatid="4817" lane="3" />
                <ENTRY entrytime="00:04:22.04" eventid="2075" heatid="4909" lane="4" />
                <ENTRY entrytime="00:09:20.58" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:20.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Niklas" gender="M" lastname="Zimmermann" nation="GER" license="345171" athleteid="2896">
              <RESULTS>
                <RESULT eventid="1763" points="507" swimtime="00:01:09.70" resultid="2897" heatid="4700" lane="5" entrytime="00:01:08.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="469" swimtime="00:00:26.06" resultid="2898" heatid="4769" lane="1" entrytime="00:00:26.26" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:31.68" eventid="1985" heatid="4844" lane="4" />
                <ENTRY entrytime="00:02:31.33" eventid="2089" heatid="4927" lane="4" />
                <ENTRY entrytime="00:00:28.55" eventid="2103" heatid="4941" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT comment="(Zeit: 19:29), Der 2. Schwimmer führte auf der Brust-Teilstrecke mehr als einen Delphin-Kick aus." eventid="2048" status="DSQ" swimtime="00:01:48.30" resultid="2902" heatid="4806" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="100" swimtime="00:00:58.45" />
                    <SPLIT distance="150" swimtime="00:01:24.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2851" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2809" number="2" reactiontime="+32" status="DSQ" />
                    <RELAYPOSITION athleteid="2846" number="3" reactiontime="+51" status="DSQ" />
                    <RELAYPOSITION athleteid="2798" number="4" reactiontime="+32" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:40.00" eventid="2232" heatid="4812" lane="1" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="2062" points="599" swimtime="00:02:03.36" resultid="2904" heatid="4807" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:37.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2786" number="1" />
                    <RELAYPOSITION athleteid="2813" number="2" />
                    <RELAYPOSITION athleteid="2794" number="3" />
                    <RELAYPOSITION athleteid="2870" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:55.00" eventid="2224" heatid="4810" lane="5" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4420" nation="GER" region="02" clubid="3434" name="TSV Neuburg">
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Fabian" gender="M" lastname="Rieß" nation="GER" license="363828" athleteid="3440">
              <RESULTS>
                <RESULT eventid="1778" points="556" swimtime="00:00:58.90" resultid="3441" heatid="4714" lane="1" entrytime="00:00:59.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="543" swimtime="00:00:27.22" resultid="3442" heatid="4741" lane="4" entrytime="00:00:27.60" />
                <RESULT eventid="1848" points="498" swimtime="00:02:13.18" resultid="3443" heatid="4789" lane="1" entrytime="00:02:15.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="150" swimtime="00:01:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1912" points="576" swimtime="00:00:26.70" resultid="5406" heatid="4744" lane="4" entrytime="00:00:27.22" />
                <RESULT eventid="1898" points="570" swimtime="00:00:58.41" resultid="5460" heatid="5465" lane="4" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:54.19" eventid="1971" heatid="4824" lane="1" />
                <ENTRY entrytime="00:01:00.26" eventid="2013" heatid="4873" lane="2" />
                <ENTRY entrytime="00:00:26.43" eventid="2103" heatid="4945" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Christina" gender="F" lastname="Wenger" nation="GER" license="162995" athleteid="3435">
              <RESULTS>
                <RESULT eventid="1756" points="573" swimtime="00:00:34.66" resultid="3436" heatid="4692" lane="1" entrytime="00:00:34.77" />
                <RESULT eventid="1799" points="495" swimtime="00:01:11.63" resultid="3437" heatid="4733" lane="5" entrytime="00:01:12.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1855" points="479" swimtime="00:00:31.15" resultid="3438" heatid="4797" lane="5" entrytime="00:00:31.05" />
                <RESULT eventid="1877" points="551" swimtime="00:00:35.12" resultid="5354" heatid="5355" lane="6" entrytime="00:00:34.66" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:01:16.16" eventid="1992" heatid="4855" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4492" nation="GER" region="02" clubid="3786" name="TSV Vaterstetten">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Christian" gender="M" lastname="Arzberger" nation="GER" license="290446" athleteid="3785">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.80" eventid="1985" heatid="4840" lane="2" />
                <ENTRY entrytime="00:02:42.51" eventid="2089" heatid="4925" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Pauline" gender="F" lastname="Breitner" nation="GER" license="273792" athleteid="3789">
              <ENTRIES>
                <ENTRY entrytime="00:02:20.01" eventid="1978" heatid="4830" lane="4" />
                <ENTRY entrytime="00:01:20.60" eventid="1992" heatid="4851" lane="5" />
                <ENTRY entrytime="00:02:40.29" eventid="2055" heatid="4896" lane="1" />
                <ENTRY entrytime="00:00:29.54" eventid="2082" heatid="4914" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Valerie" gender="F" lastname="Wende" nation="GER" license="325391" athleteid="3794">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.65" eventid="2082" heatid="4914" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5107" nation="GER" region="02" clubid="2650" name="TV 1860 Immenstadt">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Marcus" gender="M" lastname="Joas" nation="GER" license="161806" athleteid="2651">
              <RESULTS>
                <RESULT eventid="1749" points="510" swimtime="00:02:04.31" resultid="2652" heatid="4679" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="100" swimtime="00:01:00.56" />
                    <SPLIT distance="150" swimtime="00:01:32.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="464" swimtime="00:02:21.54" resultid="2653" heatid="4751" lane="5" entrytime="00:02:22.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:01:05.37" />
                    <SPLIT distance="150" swimtime="00:01:48.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="374" swimtime="00:02:26.52" resultid="2654" heatid="4787" lane="1" entrytime="00:02:21.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:11.03" />
                    <SPLIT distance="150" swimtime="00:01:48.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:58.10" eventid="1971" heatid="4815" lane="4" />
                <ENTRY entrytime="00:02:21.10" eventid="2041" heatid="4891" lane="4" />
                <ENTRY entrytime="00:04:22.25" eventid="2075" heatid="4909" lane="5" />
                <ENTRY entrytime="00:08:58.39" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:08:58.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Simon" gender="M" lastname="Joas" nation="GER" license="282570" athleteid="2659">
              <RESULTS>
                <RESULT eventid="1749" points="459" swimtime="00:02:08.80" resultid="2660" heatid="4677" lane="2" entrytime="00:02:09.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:02.22" />
                    <SPLIT distance="150" swimtime="00:01:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1834" points="423" swimtime="00:00:26.98" resultid="2661" heatid="4766" lane="5" entrytime="00:00:27.34" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:59.59" eventid="1971" heatid="4814" lane="5" />
                <ENTRY entrytime="00:04:34.09" eventid="2075" heatid="4907" lane="3" />
                <ENTRY entrytime="00:09:23.29" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:23.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4530" nation="GER" region="02" clubid="2495" name="TV 1862 Passau">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Luisa" gender="F" lastname="Roderweis" nation="GER" license="245436" athleteid="2496">
              <RESULTS>
                <RESULT eventid="1785" points="562" swimtime="00:01:06.65" resultid="2497" heatid="4724" lane="1" entrytime="00:01:06.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1813" points="542" swimtime="00:02:26.69" resultid="2498" heatid="4745" lane="4" entrytime="00:02:23.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                    <SPLIT distance="150" swimtime="00:01:49.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1827" points="684" swimtime="00:04:26.06" resultid="2499" heatid="4764" lane="5" entrytime="00:04:25.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:03.97" />
                    <SPLIT distance="150" swimtime="00:01:38.25" />
                    <SPLIT distance="200" swimtime="00:02:12.36" />
                    <SPLIT distance="250" swimtime="00:02:46.45" />
                    <SPLIT distance="300" swimtime="00:03:20.74" />
                    <SPLIT distance="350" swimtime="00:03:54.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1891" points="548" swimtime="00:01:07.24" resultid="5388" heatid="5391" lane="5" entrytime="00:01:06.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1933" points="569" swimtime="00:02:24.33" resultid="5423" heatid="4748" lane="6" entrytime="00:02:26.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:08.54" />
                    <SPLIT distance="150" swimtime="00:01:47.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:07.47" eventid="1978" heatid="4838" lane="2" />
                <ENTRY entrytime="00:09:19.00" eventid="2020" heatid="4876" lane="5">
                  <MEETINFO qualificationtime="00:09:18.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.32" eventid="2096" heatid="4936" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6812" nation="GER" region="02" clubid="2411" name="TV Kempten">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Jannes" gender="M" lastname="Schnitzer" nation="GER" license="294908" athleteid="2412">
              <RESULTS>
                <RESULT eventid="1763" points="525" swimtime="00:01:08.90" resultid="2413" heatid="4700" lane="6" entrytime="00:01:09.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="529" swimtime="00:00:59.88" resultid="2414" heatid="4713" lane="5" entrytime="00:01:00.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1820" points="568" swimtime="00:02:12.34" resultid="2415" heatid="4753" lane="6" entrytime="00:02:16.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                    <SPLIT distance="100" swimtime="00:01:01.84" />
                    <SPLIT distance="150" swimtime="00:01:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1848" points="473" swimtime="00:02:15.55" resultid="2416" heatid="4788" lane="2" entrytime="00:02:18.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="150" swimtime="00:01:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1961" points="518" swimtime="00:02:11.52" resultid="5499" heatid="5504" lane="4" entrytime="00:02:15.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                    <SPLIT distance="150" swimtime="00:01:38.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:32.53" eventid="1985" heatid="4843" lane="1" />
                <ENTRY entrytime="00:01:00.67" eventid="2013" heatid="4872" lane="2" />
                <ENTRY entrytime="00:01:03.52" eventid="2027" heatid="4879" lane="6" />
                <ENTRY entrytime="00:02:18.14" eventid="2041" heatid="4893" lane="6" />
                <ENTRY entrytime="00:02:36.99" eventid="2089" heatid="4926" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Jan" gender="M" lastname="Schuster" nation="GER" license="301516" athleteid="2422">
              <RESULTS>
                <RESULT eventid="1749" points="476" swimtime="00:02:07.20" resultid="2423" heatid="4678" lane="2" entrytime="00:02:06.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                    <SPLIT distance="100" swimtime="00:01:00.02" />
                    <SPLIT distance="150" swimtime="00:01:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1778" points="442" swimtime="00:01:03.58" resultid="2424" heatid="4711" lane="5" entrytime="00:01:02.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="385" swimtime="00:00:30.53" resultid="2425" heatid="4739" lane="5" entrytime="00:00:30.31" />
                <RESULT eventid="1834" points="492" swimtime="00:00:25.66" resultid="2426" heatid="4770" lane="3" entrytime="00:00:25.78" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:56.68" eventid="1971" heatid="4820" lane="6" />
                <ENTRY entrytime="00:01:05.05" eventid="2027" heatid="4878" lane="5" />
                <ENTRY entrytime="00:00:27.07" eventid="2103" heatid="4944" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lucas" gender="M" lastname="Willinsky" nation="GER" license="248935" athleteid="2430">
              <RESULTS>
                <RESULT eventid="1763" points="640" swimtime="00:01:04.52" resultid="2431" heatid="4701" lane="2" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1806" points="464" swimtime="00:00:28.69" resultid="2432" heatid="4741" lane="1" entrytime="00:00:28.96" />
                <RESULT eventid="1884" points="635" swimtime="00:01:04.67" resultid="5364" heatid="5368" lane="2" entrytime="00:01:04.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1912" points="482" swimtime="00:00:28.33" resultid="5416" heatid="5417" lane="6" entrytime="00:00:28.69" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:29.80" eventid="1985" heatid="4846" lane="2" />
                <ENTRY entrytime="00:01:01.14" eventid="2027" heatid="4879" lane="2" />
                <ENTRY entrytime="00:02:21.88" eventid="2089" heatid="4929" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4562" nation="GER" region="02" clubid="3230" name="TV Parsberg">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Alicia" gender="F" lastname="Urschel" nation="GER" license="300240" athleteid="3231">
              <RESULTS>
                <RESULT eventid="1059" points="564" swimtime="00:01:01.61" resultid="3232" heatid="4669" lane="4" entrytime="00:01:02.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1771" points="451" swimtime="00:05:38.29" resultid="3233" heatid="4705" lane="2" entrytime="00:05:40.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                    <SPLIT distance="150" swimtime="00:02:02.22" />
                    <SPLIT distance="200" swimtime="00:02:43.91" />
                    <SPLIT distance="250" swimtime="00:03:34.61" />
                    <SPLIT distance="300" swimtime="00:04:24.86" />
                    <SPLIT distance="350" swimtime="00:05:01.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1799" points="438" swimtime="00:01:14.61" resultid="3234" heatid="4730" lane="1" entrytime="00:01:13.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:02:18.47" eventid="1978" heatid="4831" lane="3" />
                <ENTRY entrytime="00:02:39.55" eventid="2055" heatid="4896" lane="4" />
                <ENTRY entrytime="00:00:28.43" eventid="2082" heatid="4919" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4593" nation="GER" region="02" clubid="4270" name="VfL 1860 Spfr. Bad Neustadt">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Sebastian" gender="M" lastname="Rasch" nation="GER" license="305639" athleteid="4569">
              <RESULTS>
                <RESULT eventid="1834" points="436" swimtime="00:00:26.70" resultid="4570" heatid="4768" lane="5" entrytime="00:00:26.45" />
              </RESULTS>
              <ENTRIES>
                <ENTRY entrytime="00:00:57.94" eventid="1971" heatid="4816" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1062" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="15" agemin="-1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:25.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:24.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:43.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.20">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:28.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:16.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:16.90">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1064" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="15" agemin="-1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:38.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:37.60">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:58.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:21.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:59.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:14.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.90">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:41.50">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1066" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:25.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:24.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:43.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.20">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:28.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:16.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:16.90">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1068" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:37.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.20">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:56.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:55.20">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:39.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:21.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:38.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:14.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1078" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="18" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:22.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:21.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:38.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:07.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:31.70">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:23.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:09.10">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1080" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="18" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:32.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:32.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:51.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:49.70">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:19.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:31.80">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1070" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="19" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:18.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:33.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:04.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:25.10">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:01.80">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:01.40">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:04.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1072" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="19" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:32.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:32.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:51.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:49.70">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:19.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:31.80">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="2070" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn Staffel" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:47.50">
          <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="2072" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn Staffel" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
