<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SG Fürth" version="11.61084">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Fürth" name="43. Fürther Kinderschwimmen" course="SCM" deadline="2018-11-04" hostclub="SG Fürth" hostclub.url="http://www.sgfuerth.de" organizer="SG Fürth" organizer.url="http://www.sgfuerth.de" reservecount="2" startmethod="1" timing="AUTOMATIC" state="BY" nation="GER">
      <AGEDATE value="2019-11-09" type="YEAR" />
      <POOL name="Hallebad am Scherbsgraben" lanemin="1" lanemax="6" />
      <FACILITY city="Fürth" name="Hallebad am Scherbsgraben" nation="GER" state="BY" street="Scherbsgraben 15" zip="90765" />
      <POINTTABLE pointtableid="3011" name="FINA Point Scoring" version="2018" />
      <CONTACT city="Fürth" email="meldungen@sgfuerth.de" name="Matthias Fuchs" phone="09118101172" street="Lavendelweg 47" zip="90768" />
      <SESSIONS>
        <SESSION date="2019-11-09" daytime="08:30" endtime="11:27" number="1" officialmeeting="08:15" teamleadermeeting="08:15" warmupfrom="08:00" warmupuntil="08:45">
          <EVENTS>
            <EVENT eventid="5668" gender="M" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="103" name="25m Rückenbeine ohne Brett" stroke="UNKNOWN" code="25 Rub" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7651" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7652" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7653" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7654" agemax="7" agemin="7" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7691" gender="M" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="501" name="25m Kraulbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7692" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7693" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7694" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7695" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24819" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24820" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5678" gender="M" number="5" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7659" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7660" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7661" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7662" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24812" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24813" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24814" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7696" gender="F" number="8" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="501" name="25m Kraulbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7697" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7698" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7699" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7700" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24821" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24822" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24823" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7706" gender="F" number="14" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="502" name="25m Delphinbeine o. Brett" stroke="UNKNOWN" code="25 Dob" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7707" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7708" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7709" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7710" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24835" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5674" gender="F" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="103" name="25m Rückenbeine ohne Brett" stroke="UNKNOWN" code="25 Rub" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7655" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7656" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7657" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7658" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24811" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5686" gender="M" number="9" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="101" name="25m Brustbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7667" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7668" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7669" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7670" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24824" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24825" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24826" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5664" gender="F" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7647" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7648" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7649" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7650" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24808" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24809" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24810" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5682" gender="F" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7663" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7664" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7665" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7666" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24815" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24816" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24817" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24818" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5694" gender="M" number="11" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7675" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7676" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7677" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7678" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24829" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24830" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5690" gender="F" number="10" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="101" name="25m Brustbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7671" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7672" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7673" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7674" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24827" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24828" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5698" gender="F" number="12" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7679" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7680" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7681" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7682" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24831" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24832" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24833" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1053" gender="M" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7646" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="1055" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="1054" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="2915" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24805" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24806" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24807" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7701" gender="M" number="13" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="502" name="25m Delphinbeine o. Brett" stroke="UNKNOWN" code="25 Dob" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7702" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7703" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7704" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7705" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24834" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-11-09" daytime="12:00" number="2" officialmeeting="11:30" teamleadermeeting="11:30" warmupfrom="11:00" warmupuntil="11:55">
          <EVENTS>
            <EVENT eventid="7773" gender="M" number="27" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7781" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7782" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7783" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7784" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7785" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7786" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7787" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24907" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24908" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24909" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24910" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5744" gender="F" number="26" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23817" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23818" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23819" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23820" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23821" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23822" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23823" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24898" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24899" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24900" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24901" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24902" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24903" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24904" number="7" order="7" status="SEEDED" />
                <HEAT heatid="24905" number="8" order="8" status="SEEDED" />
                <HEAT heatid="24906" number="9" order="9" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7809" gender="F" number="30" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7818" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7819" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7820" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7821" agemax="11" agemin="11" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24919" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24920" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" gender="M" number="19" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7721" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1105" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1104" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1107" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1106" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1109" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24860" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24861" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7788" gender="F" number="28" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7789" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7790" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7791" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7792" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7793" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7794" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7795" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24911" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24912" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24913" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24914" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24915" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24916" number="6" order="6" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" gender="F" number="34" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7837" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7838" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7839" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7840" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7841" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7842" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7843" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24931" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24932" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5702" gender="M" number="17" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23782" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23783" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23784" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23785" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23786" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23787" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23788" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24846" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24847" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24848" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24849" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24850" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24851" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24852" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5655" gender="M" number="37" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7870" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7871" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7872" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7873" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7874" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7875" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24946" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24947" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1177" gender="M" number="15" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7746" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7747" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7748" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7749" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7750" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7751" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24836" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24837" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24838" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5724" gender="M" number="21" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23796" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23797" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23798" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23799" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23800" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23801" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23802" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24864" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24865" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24866" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24867" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24868" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24869" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24870" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" gender="F" number="36" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7863" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7864" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7865" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7866" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7867" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7868" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7869" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24939" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24940" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24941" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24942" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24943" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24944" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24945" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5740" gender="M" number="25" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23810" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23811" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23812" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23813" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23814" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23815" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23816" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24889" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24890" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24891" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24892" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24893" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24894" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24895" number="7" order="7" status="SEEDED" />
                <HEAT heatid="24896" number="8" order="8" status="SEEDED" />
                <HEAT heatid="24897" number="9" order="9" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5661" gender="F" number="38" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7876" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7877" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7878" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7879" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7880" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7881" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24948" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7804" gender="M" number="29" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7814" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7815" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7816" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7817" agemax="11" agemin="11" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24917" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24918" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5712" gender="F" number="18" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23789" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23790" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23791" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23792" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23793" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23794" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23795" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24853" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24854" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24855" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24856" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24857" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24858" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24859" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" gender="M" number="23" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7759" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7760" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7761" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7762" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7763" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7764" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7765" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24878" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24879" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24880" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24881" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5728" gender="F" number="22" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23803" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23804" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23805" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23806" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23807" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23808" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23809" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24871" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24872" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24873" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24874" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24875" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24876" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24877" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" gender="F" number="16" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7753" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7754" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7755" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7756" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7757" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7758" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24839" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24840" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24841" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24842" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24843" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24844" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24845" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1189" gender="M" number="35" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7856" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7857" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7858" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7859" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7860" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7861" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7862" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24933" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24934" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24935" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24936" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24937" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24938" number="6" order="6" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" gender="F" number="20" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7722" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1112" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1113" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1114" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1115" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1116" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24862" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24863" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" gender="F" number="24" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7766" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7767" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7768" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7769" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7770" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7771" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7772" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24882" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24883" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24884" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24885" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24886" number="5" order="5" status="SEEDED" />
                <HEAT heatid="24887" number="6" order="6" status="SEEDED" />
                <HEAT heatid="24888" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" gender="M" number="33" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7830" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7831" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7832" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7833" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7834" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7835" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7836" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24929" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24930" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" gender="M" number="31" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23824" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23825" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23826" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23827" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23828" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23829" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23830" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24921" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24922" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24923" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1123" gender="F" number="32" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23831" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23832" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23833" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23834" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23835" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23836" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23837" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="24924" number="1" order="1" status="SEEDED" />
                <HEAT heatid="24925" number="2" order="2" status="SEEDED" />
                <HEAT heatid="24926" number="3" order="3" status="SEEDED" />
                <HEAT heatid="24927" number="4" order="4" status="SEEDED" />
                <HEAT heatid="24928" number="5" order="5" status="SEEDED" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="4224" nation="GER" region="02" clubid="23845" name="Delphin 77 Herzogenaurach">
          <ATHLETES>
            <ATHLETE birthdate="2007-01-01" firstname="Fiona" gender="F" lastname="Baumann" nation="GER" license="403954" athleteid="23846">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.62" eventid="5712" heatid="24857" lane="1" />
                <ENTRY entrytime="00:00:49.42" eventid="5728" heatid="24876" lane="6" />
                <ENTRY entrytime="00:00:39.17" eventid="5744" heatid="24905" lane="6" />
                <ENTRY entrytime="00:01:44.65" eventid="7788" heatid="24915" lane="6" />
                <ENTRY entrytime="00:00:49.02" eventid="1123" heatid="24927" lane="2" />
                <ENTRY entrytime="00:01:27.66" eventid="1195" heatid="24944" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Amelie" gender="F" lastname="Bierlmeier" nation="GER" license="426838" athleteid="23853">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.13" eventid="5712" heatid="24856" lane="3" />
                <ENTRY entrytime="00:01:01.51" eventid="5728" heatid="24873" lane="2" />
                <ENTRY entrytime="00:00:55.21" eventid="5744" heatid="24900" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lena" gender="F" lastname="Bohrer" nation="GER" license="403950" athleteid="23857">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.35" eventid="5712" heatid="24858" lane="1" />
                <ENTRY entrytime="00:00:58.95" eventid="5728" heatid="24874" lane="3" />
                <ENTRY entrytime="00:01:58.13" eventid="1135" heatid="24885" lane="4" />
                <ENTRY entrytime="00:00:48.74" eventid="5744" heatid="24902" lane="1" />
                <ENTRY entrytime="00:00:58.76" eventid="1123" heatid="24925" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Theresa" gender="F" lastname="Dellermann" nation="GER" license="410601" athleteid="23863">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.06" eventid="5712" heatid="24859" lane="5" />
                <ENTRY entrytime="00:00:44.30" eventid="5728" heatid="24877" lane="5" />
                <ENTRY entrytime="00:01:43.26" eventid="1135" heatid="24888" lane="6" />
                <ENTRY entrytime="00:00:43.23" eventid="5744" heatid="24903" lane="5" />
                <ENTRY entrytime="00:01:45.00" eventid="7788" heatid="24914" lane="4" />
                <ENTRY entrytime="00:01:10.00" eventid="1123" heatid="24924" lane="2" />
                <ENTRY entrytime="00:01:28.36" eventid="1195" heatid="24943" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Andrea Jasmin" gender="F" lastname="Erm" nation="GER" license="999999" athleteid="23871">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5712" heatid="24855" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="24874" lane="2" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="24900" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lene" gender="F" lastname="Friedrich" nation="GER" license="410600" athleteid="23875">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.51" eventid="5712" heatid="24859" lane="2" />
                <ENTRY entrytime="00:00:48.50" eventid="5728" heatid="24876" lane="5" />
                <ENTRY entrytime="00:00:37.49" eventid="5744" heatid="24905" lane="4" />
                <ENTRY entrytime="00:01:45.00" eventid="7788" heatid="24914" lane="3" />
                <ENTRY entrytime="00:01:28.40" eventid="1195" heatid="24943" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Thomas" gender="M" lastname="Hahn" nation="GER" license="999999" athleteid="23881">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5724" heatid="24864" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="24891" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Philipp" gender="M" lastname="Hardt" nation="GER" license="417042" athleteid="23884">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.19" eventid="5702" heatid="24852" lane="2" />
                <ENTRY entrytime="00:01:46.06" eventid="1141" heatid="24881" lane="1" />
                <ENTRY entrytime="00:00:37.04" eventid="5740" heatid="24896" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Simon" gender="M" lastname="Kamenik" nation="GER" license="410599" athleteid="23888">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.97" eventid="5702" heatid="24851" lane="3" />
                <ENTRY entrytime="00:00:46.40" eventid="5740" heatid="24893" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Mateo" gender="M" lastname="Kaufmair" nation="GER" license="382063" athleteid="23891">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.93" eventid="5702" heatid="24851" lane="5" />
                <ENTRY entrytime="00:00:49.19" eventid="5724" heatid="24869" lane="1" />
                <ENTRY entrytime="00:00:40.74" eventid="5740" heatid="24895" lane="5" />
                <ENTRY entrytime="00:01:44.28" eventid="7773" heatid="24909" lane="6" />
                <ENTRY entrytime="00:00:52.51" eventid="1117" heatid="24922" lane="5" />
                <ENTRY entrytime="00:01:27.37" eventid="1189" heatid="24937" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Luci" gender="F" lastname="Kitschke" nation="GER" license="417040" athleteid="23898">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.06" eventid="5712" heatid="24858" lane="5" />
                <ENTRY entrytime="00:00:50.72" eventid="5728" heatid="24875" lane="4" />
                <ENTRY entrytime="00:00:41.04" eventid="5744" heatid="24903" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Wilhelm" gender="M" lastname="Ruß" nation="GER" license="046841" athleteid="23902">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.81" eventid="5702" heatid="24850" lane="3" />
                <ENTRY entrytime="00:00:54.22" eventid="5724" heatid="24868" lane="1" />
                <ENTRY entrytime="00:01:57.00" eventid="1141" heatid="24880" lane="5" />
                <ENTRY entrytime="00:00:43.48" eventid="5740" heatid="24894" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="David" gender="M" lastname="Seefried" nation="GER" license="403947" athleteid="23907">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.67" eventid="5702" heatid="24851" lane="6" />
                <ENTRY entrytime="00:00:57.81" eventid="5724" heatid="24867" lane="1" />
                <ENTRY entrytime="00:00:45.34" eventid="5740" heatid="24893" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Jonathan" gender="M" lastname="Sopp" nation="GER" license="410602" athleteid="23911">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.51" eventid="5702" heatid="24849" lane="4" />
                <ENTRY entrytime="00:00:56.83" eventid="5724" heatid="24867" lane="2" />
                <ENTRY entrytime="00:01:57.00" eventid="1141" heatid="24880" lane="2" />
                <ENTRY entrytime="00:00:44.14" eventid="5740" heatid="24894" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emilja" gender="F" lastname="Stukelj" nation="GER" license="999999" athleteid="23916">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5712" heatid="24855" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="24873" lane="3" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="24900" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Nilaksh Vikalp" gender="M" lastname="Yadav" nation="GER" license="046836" athleteid="23920">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="5702" heatid="24850" lane="1" />
                <ENTRY entrytime="00:00:54.85" eventid="5724" heatid="24868" lane="6" />
                <ENTRY entrytime="00:00:46.07" eventid="5740" heatid="24893" lane="2" />
                <ENTRY entrytime="00:01:37.00" eventid="1189" heatid="24936" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Paul" gender="M" lastname="Zitzmann" nation="GER" license="403945" athleteid="23925">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.86" eventid="5702" heatid="24850" lane="4" />
                <ENTRY entrytime="00:00:53.73" eventid="5724" heatid="24868" lane="2" />
                <ENTRY entrytime="00:00:41.66" eventid="5740" heatid="24895" lane="6" />
                <ENTRY entrytime="00:01:45.00" eventid="7773" heatid="24908" lane="3" />
                <ENTRY entrytime="00:01:35.24" eventid="1189" heatid="24936" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6777" nation="GER" region="02" clubid="24066" name="Schwimmclub Schwandorf">
          <ATHLETES>
            <ATHLETE birthdate="2012-01-01" firstname="Luca" gender="M" lastname="Daucher" nation="GER" license="404783" athleteid="24067">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.02" eventid="1053" heatid="24807" lane="2" />
                <ENTRY entrytime="00:00:28.82" eventid="5678" heatid="24814" lane="4" />
                <ENTRY entrytime="00:00:36.77" eventid="7691" heatid="24820" lane="4" />
                <ENTRY entrytime="00:00:31.80" eventid="5694" heatid="24830" lane="2" />
                <ENTRY entrytime="NT" eventid="7701" heatid="24834" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Carlotta" gender="F" lastname="Fleischmann" nation="GER" license="374674" athleteid="24073">
              <ENTRIES>
                <ENTRY entrytime="00:03:30.08" eventid="1183" heatid="24842" lane="5" />
                <ENTRY entrytime="00:00:49.26" eventid="5728" heatid="24876" lane="1" />
                <ENTRY entrytime="00:01:56.51" eventid="1135" heatid="24885" lane="3" />
                <ENTRY entrytime="00:01:45.08" eventid="7788" heatid="24914" lane="2" />
                <ENTRY entrytime="00:00:50.51" eventid="1123" heatid="24927" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lucie" gender="F" lastname="Gebele" nation="GER" license="405006" athleteid="24085">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.57" eventid="5712" heatid="24854" lane="4" />
                <ENTRY entrytime="00:01:15.55" eventid="5728" heatid="24871" lane="2" />
                <ENTRY entrytime="NT" eventid="1135" heatid="24882" lane="2" />
                <ENTRY entrytime="00:01:09.03" eventid="5744" heatid="24898" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Helena" gender="F" lastname="Gäntzle" nation="GER" license="405005" athleteid="24079">
              <ENTRIES>
                <ENTRY entrytime="00:03:18.57" eventid="1183" heatid="24843" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="1111" heatid="24863" lane="6" />
                <ENTRY entrytime="00:00:40.34" eventid="5744" heatid="24904" lane="1" />
                <ENTRY entrytime="00:01:44.40" eventid="7788" heatid="24915" lane="1" />
                <ENTRY entrytime="00:00:46.94" eventid="1123" heatid="24927" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Andreas" gender="M" lastname="Hiltl" nation="GER" license="371456" athleteid="24090">
              <ENTRIES>
                <ENTRY entrytime="00:04:12.62" eventid="1177" heatid="24836" lane="1" />
                <ENTRY entrytime="00:01:05.54" eventid="5702" heatid="24847" lane="4" />
                <ENTRY entrytime="00:01:00.48" eventid="5724" heatid="24866" lane="2" />
                <ENTRY entrytime="00:00:45.60" eventid="5740" heatid="24893" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Knerer" nation="GER" license="404785" athleteid="24095">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5674" heatid="24811" lane="1" />
                <ENTRY entrytime="00:00:31.86" eventid="5682" heatid="24818" lane="5" />
                <ENTRY entrytime="00:00:44.97" eventid="7696" heatid="24823" lane="1" />
                <ENTRY entrytime="00:00:36.75" eventid="5698" heatid="24833" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emma" gender="F" lastname="Köhn" nation="GER" license="418818" athleteid="24100">
              <ENTRIES>
                <ENTRY entrytime="00:03:43.16" eventid="1183" heatid="24841" lane="1" />
                <ENTRY entrytime="00:00:56.40" eventid="5712" heatid="24857" lane="4" />
                <ENTRY entrytime="00:00:42.23" eventid="5744" heatid="24903" lane="2" />
                <ENTRY entrytime="00:01:55.44" eventid="7788" heatid="24913" lane="4" />
                <ENTRY entrytime="00:00:57.29" eventid="1123" heatid="24925" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Abby" gender="F" lastname="Lukas" nation="GER" license="374673" athleteid="24106">
              <ENTRIES>
                <ENTRY entrytime="00:03:27.71" eventid="1183" heatid="24842" lane="4" />
                <ENTRY entrytime="00:02:15.00" eventid="1111" heatid="24862" lane="2" />
                <ENTRY entrytime="00:00:45.59" eventid="5744" heatid="24902" lane="3" />
                <ENTRY entrytime="00:02:01.46" eventid="7788" heatid="24913" lane="1" />
                <ENTRY entrytime="00:00:57.34" eventid="1123" heatid="24925" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Aleksei" gender="M" lastname="Malikoski" nation="GER" license="390306" athleteid="24112">
              <ENTRIES>
                <ENTRY entrytime="00:03:16.36" eventid="1177" heatid="24837" lane="1" />
                <ENTRY entrytime="00:00:49.75" eventid="5724" heatid="24869" lane="6" />
                <ENTRY entrytime="00:00:38.19" eventid="5740" heatid="24896" lane="1" />
                <ENTRY entrytime="00:00:55.24" eventid="1117" heatid="24921" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Eva" gender="F" lastname="Matthes" nation="GER" license="000000" athleteid="24117">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.41" eventid="5664" heatid="24809" lane="3" />
                <ENTRY entrytime="NT" eventid="5674" heatid="24811" lane="2" />
                <ENTRY entrytime="00:00:37.55" eventid="5682" heatid="24817" lane="4" />
                <ENTRY entrytime="00:00:34.37" eventid="5690" heatid="24828" lane="4" />
                <ENTRY entrytime="00:00:42.56" eventid="5698" heatid="24832" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Ida" gender="F" lastname="Matthes" nation="GER" license="416783" athleteid="24123">
              <ENTRIES>
                <ENTRY entrytime="00:05:46.11" eventid="1183" heatid="24839" lane="2" />
                <ENTRY entrytime="00:00:59.53" eventid="5712" heatid="24856" lane="5" />
                <ENTRY entrytime="00:02:16.28" eventid="1135" heatid="24883" lane="2" />
                <ENTRY entrytime="00:00:54.36" eventid="5744" heatid="24901" lane="1" />
                <ENTRY entrytime="00:02:17.73" eventid="7788" heatid="24911" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Paulina" gender="F" lastname="Plößl" nation="GER" license="374754" athleteid="24129">
              <ENTRIES>
                <ENTRY entrytime="00:04:10.70" eventid="1183" heatid="24839" lane="3" />
                <ENTRY entrytime="00:00:58.52" eventid="5712" heatid="24856" lane="4" />
                <ENTRY entrytime="00:02:06.48" eventid="1135" heatid="24884" lane="1" />
                <ENTRY entrytime="00:02:16.88" eventid="7788" heatid="24911" lane="2" />
                <ENTRY entrytime="00:00:59.17" eventid="1123" heatid="24924" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Hanna" gender="F" lastname="Rieder" nation="GER" license="390308" athleteid="24135">
              <ENTRIES>
                <ENTRY entrytime="00:03:39.57" eventid="1183" heatid="24841" lane="2" />
                <ENTRY entrytime="00:02:20.00" eventid="1111" heatid="24862" lane="5" />
                <ENTRY entrytime="00:00:46.31" eventid="5744" heatid="24902" lane="4" />
                <ENTRY entrytime="00:02:02.10" eventid="7788" heatid="24913" lane="6" />
                <ENTRY entrytime="00:00:56.68" eventid="1123" heatid="24925" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Victoria" gender="F" lastname="Schmid" nation="GER" license="421993" athleteid="24141">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.75" eventid="5728" heatid="24871" lane="5" />
                <ENTRY entrytime="00:01:10.29" eventid="5744" heatid="24898" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leonie" gender="F" lastname="Seger" nation="GER" license="390311" athleteid="24144">
              <ENTRIES>
                <ENTRY entrytime="00:03:18.65" eventid="1183" heatid="24843" lane="4" />
                <ENTRY entrytime="00:00:50.16" eventid="5728" heatid="24875" lane="3" />
                <ENTRY entrytime="00:00:40.11" eventid="5744" heatid="24904" lane="2" />
                <ENTRY entrytime="00:01:50.08" eventid="7788" heatid="24914" lane="5" />
                <ENTRY entrytime="00:00:50.68" eventid="1123" heatid="24926" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Zoe" gender="F" lastname="Seger" nation="GER" license="390312" athleteid="24150">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.30" eventid="5712" heatid="24858" lane="2" />
                <ENTRY entrytime="00:02:05.00" eventid="1135" heatid="24884" lane="2" />
                <ENTRY entrytime="00:00:43.25" eventid="5744" heatid="24903" lane="1" />
                <ENTRY entrytime="00:02:05.36" eventid="7788" heatid="24912" lane="2" />
                <ENTRY entrytime="00:00:48.60" eventid="1123" heatid="24927" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Anton" gender="M" lastname="Stiegler" nation="GER" license="421391" athleteid="24156">
              <ENTRIES>
                <ENTRY entrytime="00:01:22.69" eventid="5702" heatid="24846" lane="2" />
                <ENTRY entrytime="00:01:31.33" eventid="5724" heatid="24864" lane="2" />
                <ENTRY entrytime="00:01:38.51" eventid="5740" heatid="24889" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lara" gender="F" lastname="Wachtel" nation="GER" license="404786" athleteid="24160">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.50" eventid="5664" heatid="24810" lane="3" />
                <ENTRY entrytime="00:00:26.22" eventid="5682" heatid="24818" lane="4" />
                <ENTRY entrytime="00:00:47.95" eventid="5690" heatid="24828" lane="6" />
                <ENTRY entrytime="00:00:31.11" eventid="5698" heatid="24833" lane="4" />
                <ENTRY entrytime="NT" eventid="7706" heatid="24835" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Pauline" gender="F" lastname="Wiederer" nation="GER" license="390242" athleteid="24166">
              <ENTRIES>
                <ENTRY entrytime="00:03:53.12" eventid="1183" heatid="24840" lane="4" />
                <ENTRY entrytime="00:00:48.28" eventid="5728" heatid="24876" lane="2" />
                <ENTRY entrytime="00:02:05.54" eventid="1135" heatid="24884" lane="5" />
                <ENTRY entrytime="00:02:01.33" eventid="7788" heatid="24913" lane="5" />
                <ENTRY entrytime="00:00:54.49" eventid="1123" heatid="24926" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lina-Marie" gender="F" lastname="Zimmermann-Grünauer" nation="GER" license="420366" athleteid="24172">
              <ENTRIES>
                <ENTRY entrytime="00:04:11.21" eventid="1183" heatid="24839" lane="4" />
                <ENTRY entrytime="00:01:00.73" eventid="5712" heatid="24856" lane="6" />
                <ENTRY entrytime="00:02:10.32" eventid="1135" heatid="24883" lane="4" />
                <ENTRY entrytime="00:02:10.80" eventid="7788" heatid="24911" lane="3" />
                <ENTRY entrytime="00:01:03.81" eventid="1123" heatid="24924" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4302" nation="GER" region="02" clubid="24664" name="Schwimmfreunde Pegnitz">
          <ATHLETES>
            <ATHLETE birthdate="2008-01-01" firstname="Max" gender="M" lastname="Appelhans" nation="GER" license="382234" athleteid="24665">
              <ENTRIES>
                <ENTRY entrytime="00:03:16.75" eventid="1177" heatid="24837" lane="6" />
                <ENTRY entrytime="00:00:46.63" eventid="5724" heatid="24870" lane="6" />
                <ENTRY entrytime="00:00:38.77" eventid="5740" heatid="24895" lane="3" />
                <ENTRY entrytime="00:00:50.73" eventid="1117" heatid="24922" lane="2" />
                <ENTRY entrytime="00:01:29.14" eventid="1189" heatid="24937" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Hanna" gender="F" lastname="Büttner" nation="GER" license="419941" athleteid="24671">
              <ENTRIES>
                <ENTRY entrytime="00:03:30.45" eventid="1183" heatid="24842" lane="1" />
                <ENTRY entrytime="00:00:40.73" eventid="5728" heatid="24877" lane="4" />
                <ENTRY entrytime="00:01:31.23" eventid="1171" heatid="24932" lane="4" />
                <ENTRY entrytime="00:03:29.29" eventid="5661" heatid="24948" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jan" gender="M" lastname="Büttner" nation="GER" license="419943" athleteid="24676">
              <ENTRIES>
                <ENTRY entrytime="00:03:32.96" eventid="1177" heatid="24836" lane="3" />
                <ENTRY entrytime="00:00:46.80" eventid="5724" heatid="24869" lane="4" />
                <ENTRY entrytime="00:00:40.45" eventid="5740" heatid="24895" lane="2" />
                <ENTRY entrytime="00:01:48.00" eventid="7773" heatid="24908" lane="4" />
                <ENTRY entrytime="00:01:32.17" eventid="1189" heatid="24936" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Annika" gender="F" lastname="Reichel" nation="GER" license="419942" athleteid="24682">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.00" eventid="1183" heatid="24844" lane="2" />
                <ENTRY entrytime="00:00:46.65" eventid="5712" heatid="24859" lane="4" />
                <ENTRY entrytime="00:01:39.93" eventid="1135" heatid="24888" lane="5" />
                <ENTRY entrytime="00:03:29.82" eventid="5661" heatid="24948" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5147" nation="GER" region="02" clubid="23839" name="Schwimmgemeinschaft Fürth">
          <ATHLETES>
            <ATHLETE birthdate="2007-12-08" firstname="Philipp" gender="M" lastname="Adler" nation="GER" license="407267" athleteid="23977">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.87" entrycourse="SCM" eventid="5702" heatid="24848" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="7773" heatid="24907" lane="5" />
                <ENTRY entrytime="00:01:56.04" entrycourse="SCM" eventid="1189" heatid="24934" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Aidan" gender="M" lastname="Amelong" nation="GER" license="370804" athleteid="24492">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.74" eventid="5702" heatid="24851" lane="4" />
                <ENTRY entrytime="00:01:45.72" eventid="1141" heatid="24881" lane="5" />
                <ENTRY entrytime="00:01:18.54" eventid="1189" heatid="24937" lane="4" />
                <ENTRY entrytime="00:01:36.73" eventid="7773" heatid="24909" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Sina" gender="F" lastname="Amelong" nation="GER" license="378026" athleteid="24687">
              <ENTRIES>
                <ENTRY entrytime="00:03:23.58" eventid="1183" heatid="24843" lane="1" />
                <ENTRY entrytime="00:02:00.00" eventid="1111" heatid="24862" lane="3" />
                <ENTRY entrytime="00:01:05.80" eventid="7788" heatid="24916" lane="3" />
                <ENTRY entrytime="00:01:30.19" eventid="1195" heatid="24943" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sinan" gender="M" lastname="Arpert" nation="GER" license="297748" athleteid="24497">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.13" eventid="5702" heatid="24852" lane="3" />
                <ENTRY entrytime="00:01:27.19" eventid="1141" heatid="24881" lane="4" />
                <ENTRY entrytime="00:01:27.46" eventid="7773" heatid="24910" lane="2" />
                <ENTRY entrytime="00:03:02.69" eventid="5655" heatid="24947" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-03-07" firstname="Daniel" gender="M" lastname="Asev-Ajiyev" nation="GER" license="356304" athleteid="23981">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.81" entrycourse="SCM" eventid="5702" heatid="24850" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.35" entrycourse="SCM" eventid="5724" heatid="24867" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.82" entrycourse="SCM" eventid="5740" heatid="24894" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Marie" gender="F" lastname="Auerbach" nation="GER" license="391816" athleteid="24502">
              <ENTRIES>
                <ENTRY entrytime="00:01:47.35" eventid="1111" heatid="24863" lane="5" />
                <ENTRY entrytime="00:01:48.99" eventid="1135" heatid="24887" lane="5" />
                <ENTRY entrytime="00:01:39.94" eventid="7788" heatid="24915" lane="5" />
                <ENTRY entrytime="00:00:46.47" eventid="1123" heatid="24928" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lara" gender="F" lastname="Bamberger" nation="GER" license="362930" athleteid="24178">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.86" eventid="5712" heatid="24858" lane="4" />
                <ENTRY entrytime="00:00:47.65" eventid="5728" heatid="24876" lane="3" />
                <ENTRY entrytime="00:00:38.11" eventid="5744" heatid="24905" lane="2" />
                <ENTRY entrytime="00:00:50.74" eventid="1123" heatid="24926" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-23" firstname="Rebekka" gender="F" lastname="Behring" nation="GER" license="407272" athleteid="24482">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.00" eventid="5728" heatid="24873" lane="5" />
                <ENTRY entrytime="00:01:04.00" eventid="5744" heatid="24899" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Max Eric" gender="M" lastname="Besecke" nation="GER" license="406834" athleteid="24692">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1141" heatid="24879" lane="3" />
                <ENTRY entrytime="00:01:02.37" eventid="5740" heatid="24891" lane="6" />
                <ENTRY entrytime="00:02:05.00" eventid="1189" heatid="24934" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Alarice" gender="F" lastname="Bitz" nation="GER" athleteid="24696">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="24808" lane="6" />
                <ENTRY entrytime="NT" eventid="5682" heatid="24815" lane="5" />
                <ENTRY entrytime="NT" eventid="5690" heatid="24827" lane="6" />
                <ENTRY entrytime="NT" eventid="5698" heatid="24831" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Benedek" gender="M" lastname="Boha" nation="GER" license="666666" athleteid="24701">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1177" heatid="24836" lane="6" />
                <ENTRY entrytime="00:01:50.00" eventid="1141" heatid="24880" lane="4" />
                <ENTRY entrytime="NT" eventid="7773" heatid="24907" lane="1" />
                <ENTRY entrytime="00:01:40.00" eventid="1189" heatid="24936" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Dina" gender="F" lastname="Boha" nation="GER" license="391813" athleteid="24507">
              <ENTRIES>
                <ENTRY entrytime="00:02:47.51" eventid="1183" heatid="24845" lane="3" />
                <ENTRY entrytime="00:01:38.74" eventid="1135" heatid="24888" lane="2" />
                <ENTRY entrytime="00:01:30.09" eventid="7788" heatid="24916" lane="2" />
                <ENTRY entrytime="00:01:13.15" eventid="1195" heatid="24945" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-04-17" firstname="Daniel" gender="M" lastname="Bramigk" nation="GER" license="420770" athleteid="23990">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.48" entrycourse="SCM" eventid="5724" heatid="24867" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:48.64" entrycourse="SCM" eventid="5740" heatid="24893" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:44.78" entrycourse="LCM" eventid="1189" heatid="24935" lane="2">
                  <MEETINFO course="LCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Anastasia" gender="F" lastname="Chochlow" nation="GER" license="392745" athleteid="24706">
              <ENTRIES>
                <ENTRY entrytime="00:03:29.58" eventid="1183" heatid="24842" lane="2" />
                <ENTRY entrytime="00:00:02.00" eventid="1111" heatid="24863" lane="3" />
                <ENTRY entrytime="00:01:53.07" eventid="7788" heatid="24914" lane="6" />
                <ENTRY entrytime="00:01:35.19" eventid="1195" heatid="24942" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lena" gender="F" lastname="Clausen" nation="GER" license="420945" athleteid="24512">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.53" eventid="5712" heatid="24855" lane="2" />
                <ENTRY entrytime="00:01:04.27" eventid="5728" heatid="24872" lane="3" />
                <ENTRY entrytime="00:01:01.92" eventid="5744" heatid="24899" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="7809" heatid="24919" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Simon" gender="M" lastname="Clausen" nation="GER" athleteid="24517">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.38" eventid="1053" heatid="24806" lane="2" />
                <ENTRY entrytime="00:00:50.00" eventid="7691" heatid="24820" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5686" heatid="24825" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Simon" gender="M" lastname="Dieret" nation="GER" license="331161" athleteid="23840">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.62" eventid="5724" heatid="24870" lane="5" />
                <ENTRY entrytime="00:00:35.24" eventid="5740" heatid="24897" lane="6" />
                <ENTRY entrytime="00:01:33.75" eventid="7773" heatid="24909" lane="3" />
                <ENTRY entrytime="00:00:41.54" eventid="1117" heatid="24923" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Daniel" gender="M" lastname="Ehnis" nation="GER" license="378024" athleteid="24711">
              <ENTRIES>
                <ENTRY entrytime="00:03:57.93" eventid="1177" heatid="24836" lane="2" />
                <ENTRY entrytime="00:02:03.30" eventid="1141" heatid="24880" lane="6" />
                <ENTRY entrytime="00:02:06.48" eventid="7773" heatid="24907" lane="4" />
                <ENTRY entrytime="00:01:45.32" eventid="1189" heatid="24935" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Julia" gender="F" lastname="Ehnis" nation="GER" athleteid="24716">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.36" eventid="5664" heatid="24810" lane="1" />
                <ENTRY entrytime="00:00:48.60" eventid="5682" heatid="24816" lane="3" />
                <ENTRY entrytime="00:00:48.00" eventid="7696" heatid="24823" lane="6" />
                <ENTRY entrytime="00:00:45.51" eventid="5698" heatid="24832" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-02-15" firstname="Jakob" gender="M" lastname="Freund" nation="GER" license="331165" athleteid="23994">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.37" entrycourse="SCM" eventid="5702" heatid="24850" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.97" entrycourse="SCM" eventid="5724" heatid="24866" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.92" entrycourse="SCM" eventid="5740" heatid="24892" lane="2">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.23" entrycourse="SCM" eventid="1117" heatid="24921" lane="2">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lia Sophie" gender="F" lastname="Fuchs" nation="GER" license="420938" athleteid="24721">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.38" eventid="5664" heatid="24810" lane="6" />
                <ENTRY entrytime="NT" eventid="5674" heatid="24811" lane="5" />
                <ENTRY entrytime="00:00:31.58" eventid="5682" heatid="24818" lane="2" />
                <ENTRY entrytime="00:00:33.75" eventid="5698" heatid="24833" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Linnea Emilia" gender="F" lastname="Glößinger" nation="GER" license="389377" athleteid="24726">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.84" eventid="5664" heatid="24810" lane="2" />
                <ENTRY entrytime="00:00:36.63" eventid="5682" heatid="24817" lane="3" />
                <ENTRY entrytime="00:00:00.50" eventid="5690" heatid="24828" lane="3" />
                <ENTRY entrytime="00:00:36.14" eventid="5698" heatid="24833" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Anton" gender="M" lastname="Grießinger" nation="GER" license="362946" athleteid="24521">
              <ENTRIES>
                <ENTRY entrytime="00:01:26.58" eventid="1103" heatid="24861" lane="4" />
                <ENTRY entrytime="00:01:40.44" eventid="1141" heatid="24881" lane="2" />
                <ENTRY entrytime="00:01:27.92" eventid="7773" heatid="24910" lane="1" />
                <ENTRY entrytime="00:01:12.39" eventid="1189" heatid="24938" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Annika" gender="F" lastname="Haas" nation="GER" license="555555" athleteid="24183">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="24874" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-12-18" firstname="Maximilian" gender="M" lastname="Hahn" nation="GER" license="406837" athleteid="24485">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5702" heatid="24847" lane="3" />
                <ENTRY entrytime="00:01:02.55" entrycourse="SCM" eventid="5724" heatid="24866" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-17" name="Vereinsmeisterschaft 2019" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.52" entrycourse="SCM" eventid="5740" heatid="24892" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-17" name="Vereinsmeisterschaft 2019" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lilith" gender="F" lastname="Heidenreich" nation="GER" license="420940" athleteid="24526">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.43" eventid="5712" heatid="24854" lane="2" />
                <ENTRY entrytime="00:01:05.81" eventid="5744" heatid="24899" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Louisa" gender="F" lastname="Heidenreich" nation="GER" license="420942" athleteid="24529">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.76" eventid="5664" heatid="24809" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="24831" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Luisa" gender="F" lastname="Heyert" nation="GER" license="347335" athleteid="24532">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.65" eventid="5712" heatid="24858" lane="3" />
                <ENTRY entrytime="00:00:42.56" eventid="5728" heatid="24877" lane="2" />
                <ENTRY entrytime="00:01:30.77" eventid="7788" heatid="24916" lane="1" />
                <ENTRY entrytime="00:01:20.37" eventid="1195" heatid="24945" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Tobias" gender="M" lastname="Heyert" nation="GER" license="306630" athleteid="24537">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.65" eventid="5724" heatid="24870" lane="3" />
                <ENTRY entrytime="00:00:29.85" eventid="5740" heatid="24897" lane="4" />
                <ENTRY entrytime="00:01:16.78" eventid="1165" heatid="24930" lane="3" />
                <ENTRY entrytime="00:02:49.82" eventid="5655" heatid="24947" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Alissa" gender="F" lastname="Hilz" nation="GER" athleteid="24731">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="24853" lane="4" />
                <ENTRY entrytime="NT" eventid="1135" heatid="24882" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Julianna" gender="F" lastname="Jahn" nation="GER" athleteid="24542">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5728" heatid="24872" lane="6" />
                <ENTRY entrytime="00:01:10.00" eventid="5744" heatid="24898" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Emil" gender="M" lastname="Jeske" nation="GER" license="378027" athleteid="24734">
              <ENTRIES>
                <ENTRY entrytime="00:03:02.16" eventid="1177" heatid="24837" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="1103" heatid="24860" lane="2" />
                <ENTRY entrytime="00:01:33.44" eventid="1165" heatid="24930" lane="5" />
                <ENTRY entrytime="00:03:00.00" eventid="5655" heatid="24947" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Vanessa" gender="F" lastname="Kenner" nation="GER" license="362937" athleteid="24185">
              <ENTRIES>
                <ENTRY entrytime="00:03:50.34" eventid="1183" heatid="24840" lane="3" />
                <ENTRY entrytime="00:02:00.99" eventid="1171" heatid="24931" lane="3" />
                <ENTRY entrytime="00:04:45.00" eventid="5661" heatid="24948" lane="5" />
                <ENTRY entrytime="00:02:10.00" eventid="1111" heatid="24862" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Max" gender="M" lastname="Keyser" nation="GER" license="420769" athleteid="24190">
              <ENTRIES>
                <ENTRY entrytime="00:02:59.12" eventid="1177" heatid="24837" lane="3" />
                <ENTRY entrytime="00:01:40.00" eventid="1103" heatid="24861" lane="1" />
                <ENTRY entrytime="00:03:40.00" eventid="5655" heatid="24946" lane="4" />
                <ENTRY entrytime="00:00:33.21" eventid="5740" heatid="24897" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Timm" gender="M" lastname="Laus" nation="GER" license="362943" athleteid="24195">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.69" eventid="5702" heatid="24849" lane="3" />
                <ENTRY entrytime="00:00:55.63" eventid="5724" heatid="24867" lane="4" />
                <ENTRY entrytime="00:02:00.00" eventid="7773" heatid="24908" lane="1" />
                <ENTRY entrytime="00:01:55.00" eventid="1165" heatid="24929" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Luca" gender="M" lastname="Lautenschlager" nation="GER" license="404302" athleteid="23931">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.06" eventid="1053" heatid="24807" lane="4" />
                <ENTRY entrytime="00:00:35.41" eventid="5678" heatid="24813" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="24826" lane="1" />
                <ENTRY entrytime="00:00:39.64" eventid="5694" heatid="24829" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Nils" gender="M" lastname="Lautenschlager" nation="GER" license="372637" athleteid="23936">
              <ENTRIES>
                <ENTRY entrytime="00:02:15.00" eventid="1141" heatid="24878" lane="2" />
                <ENTRY entrytime="00:00:55.19" eventid="5724" heatid="24867" lane="3" />
                <ENTRY entrytime="00:00:27.00" eventid="7804" heatid="24918" lane="2" />
                <ENTRY entrytime="00:02:15.00" eventid="1189" heatid="24933" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Edwin" gender="M" lastname="Lichtenwald" nation="GER" athleteid="24739">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.31" eventid="1053" heatid="24806" lane="4" />
                <ENTRY entrytime="00:00:33.54" eventid="5678" heatid="24814" lane="5" />
                <ENTRY entrytime="00:00:00.50" eventid="5686" heatid="24826" lane="2" />
                <ENTRY entrytime="00:00:37.22" eventid="5694" heatid="24829" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Livia" gender="F" lastname="Lichtenwald" nation="GER" license="393386" athleteid="24744">
              <ENTRIES>
                <ENTRY entrytime="00:03:22.51" eventid="1183" heatid="24843" lane="5" />
                <ENTRY entrytime="00:01:48.78" eventid="1111" heatid="24863" lane="1" />
                <ENTRY entrytime="00:01:46.72" eventid="1135" heatid="24887" lane="2" />
                <ENTRY entrytime="00:01:31.33" eventid="1195" heatid="24943" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Finn" gender="M" lastname="Martin" nation="GER" license="355301" athleteid="24200">
              <ENTRIES>
                <ENTRY entrytime="00:03:01.34" eventid="1177" heatid="24837" lane="4" />
                <ENTRY entrytime="00:01:40.91" eventid="1103" heatid="24860" lane="3" />
                <ENTRY entrytime="00:00:33.03" eventid="5740" heatid="24897" lane="2" />
                <ENTRY entrytime="00:03:45.00" eventid="5655" heatid="24946" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ida" gender="F" lastname="Martin" nation="GER" license="362939" athleteid="24205">
              <ENTRIES>
                <ENTRY entrytime="00:03:36.02" eventid="1183" heatid="24841" lane="4" />
                <ENTRY entrytime="00:02:17.91" eventid="1135" heatid="24883" lane="5" />
                <ENTRY entrytime="00:00:55.59" eventid="1123" heatid="24925" lane="3" />
                <ENTRY entrytime="00:01:42.54" eventid="1195" heatid="24941" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Cosima" gender="F" lastname="Nahr" nation="GER" license="376904" athleteid="23941">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.56" eventid="5728" heatid="24875" lane="2" />
                <ENTRY entrytime="00:01:58.57" eventid="1135" heatid="24885" lane="5" />
                <ENTRY entrytime="00:00:26.00" eventid="7809" heatid="24920" lane="4" />
                <ENTRY entrytime="00:02:10.00" eventid="1195" heatid="24939" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Julius" gender="M" lastname="Nahr" nation="GER" license="416999" athleteid="23946">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.06" eventid="1053" heatid="24806" lane="1" />
                <ENTRY entrytime="00:00:40.00" eventid="7691" heatid="24820" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="24826" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Julia" gender="F" lastname="Okner" nation="GER" athleteid="23950">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.38" eventid="5712" heatid="24853" lane="3" />
                <ENTRY entrytime="00:01:30.12" eventid="5744" heatid="24898" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jonas" gender="M" lastname="Penz" nation="GER" license="392570" athleteid="24210">
              <ENTRIES>
                <ENTRY entrytime="00:04:00.43" eventid="1177" heatid="24836" lane="5" />
                <ENTRY entrytime="00:00:53.53" eventid="5724" heatid="24868" lane="4" />
                <ENTRY entrytime="00:00:41.53" eventid="5740" heatid="24895" lane="1" />
                <ENTRY entrytime="00:01:42.69" eventid="1189" heatid="24935" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lara" gender="F" lastname="Penz" nation="GER" license="362938" athleteid="24215">
              <ENTRIES>
                <ENTRY entrytime="00:03:26.58" eventid="1183" heatid="24842" lane="3" />
                <ENTRY entrytime="00:00:36.68" eventid="5744" heatid="24906" lane="6" />
                <ENTRY entrytime="00:00:44.22" eventid="1123" heatid="24928" lane="5" />
                <ENTRY entrytime="00:03:37.69" eventid="5661" heatid="24948" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-13" firstname="Laurenz" gender="M" lastname="Raum" nation="GER" license="392567" athleteid="24489">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.00" eventid="5702" heatid="24848" lane="2" />
                <ENTRY entrytime="00:00:59.00" eventid="5740" heatid="24891" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lian" gender="M" lastname="Richter" nation="GER" license="406841" athleteid="24749">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1141" heatid="24879" lane="2" />
                <ENTRY entrytime="00:00:29.15" eventid="7804" heatid="24918" lane="5" />
                <ENTRY entrytime="NT" eventid="1165" heatid="24929" lane="2" />
                <ENTRY entrytime="00:02:25.28" eventid="1189" heatid="24933" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lisa" gender="F" lastname="Rischbeck" nation="GER" license="666666" athleteid="24754">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1135" heatid="24884" lane="4" />
                <ENTRY entrytime="NT" eventid="7788" heatid="24911" lane="1" />
                <ENTRY entrytime="NT" eventid="7809" heatid="24919" lane="1" />
                <ENTRY entrytime="00:02:00.00" eventid="1195" heatid="24940" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Theo" gender="M" lastname="Rischbeck" nation="GER" license="666666" athleteid="24759">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.19" eventid="1053" heatid="24807" lane="6" />
                <ENTRY entrytime="00:00:33.82" eventid="5678" heatid="24814" lane="1" />
                <ENTRY entrytime="00:00:00.45" eventid="5686" heatid="24826" lane="3" />
                <ENTRY entrytime="00:00:36.23" eventid="5694" heatid="24830" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ronja" gender="F" lastname="Rosenthal" nation="GER" license="389376" athleteid="24764">
              <ENTRIES>
                <ENTRY entrytime="00:03:57.10" eventid="1183" heatid="24840" lane="5" />
                <ENTRY entrytime="00:01:49.69" eventid="1135" heatid="24887" lane="6" />
                <ENTRY entrytime="00:01:39.75" eventid="1171" heatid="24932" lane="2" />
                <ENTRY entrytime="00:01:32.28" eventid="1195" heatid="24942" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Leana Isabel" gender="F" lastname="Rother" nation="GER" license="379366" athleteid="23953">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.56" eventid="5728" heatid="24875" lane="5" />
                <ENTRY entrytime="00:01:58.44" eventid="1135" heatid="24885" lane="2" />
                <ENTRY entrytime="00:00:26.00" eventid="7809" heatid="24920" lane="2" />
                <ENTRY entrytime="00:01:53.91" eventid="1195" heatid="24941" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Theo" gender="M" lastname="Rother" nation="GER" athleteid="24769">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.25" eventid="1053" heatid="24807" lane="5" />
                <ENTRY entrytime="00:00:29.52" eventid="5678" heatid="24814" lane="2" />
                <ENTRY entrytime="00:00:00.45" eventid="5686" heatid="24826" lane="4" />
                <ENTRY entrytime="00:00:31.79" eventid="5694" heatid="24830" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Timon Sebastian" gender="M" lastname="Rother" nation="GER" license="406840" athleteid="23958">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.19" eventid="1053" heatid="24807" lane="1" />
                <ENTRY entrytime="00:00:35.43" eventid="5678" heatid="24813" lane="4" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="24826" lane="6" />
                <ENTRY entrytime="00:00:36.50" eventid="5694" heatid="24829" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-10-21" firstname="Lisa" gender="F" lastname="Rutkowski" nation="GER" license="377885" athleteid="23999">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.51" entrycourse="SCM" eventid="5712" heatid="24859" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.27" entrycourse="SCM" eventid="5744" heatid="24904" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.15" entrycourse="SCM" eventid="1123" heatid="24928" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Jonathan" gender="M" lastname="Sandig" nation="GER" license="413757" athleteid="24220">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.34" eventid="5702" heatid="24852" lane="5" />
                <ENTRY entrytime="00:02:07.09" eventid="1141" heatid="24879" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="7773" heatid="24908" lane="6" />
                <ENTRY entrytime="00:01:41.74" eventid="1189" heatid="24935" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Diana" gender="F" lastname="Satsevich" nation="GER" license="391760" athleteid="24545">
              <ENTRIES>
                <ENTRY entrytime="00:02:55.25" eventid="1183" heatid="24845" lane="2" />
                <ENTRY entrytime="00:00:46.46" eventid="5728" heatid="24877" lane="6" />
                <ENTRY entrytime="00:01:35.90" eventid="7788" heatid="24915" lane="4" />
                <ENTRY entrytime="00:01:19.65" eventid="1195" heatid="24945" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Jan" gender="M" lastname="Schafner" nation="GER" license="406833" athleteid="24774">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1141" heatid="24879" lane="4" />
                <ENTRY entrytime="00:00:35.00" eventid="7804" heatid="24917" lane="4" />
                <ENTRY entrytime="NT" eventid="1165" heatid="24929" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1189" heatid="24934" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Maximilian" gender="M" lastname="Schechtel" nation="GER" athleteid="24779">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="24805" lane="2" />
                <ENTRY entrytime="NT" eventid="5678" heatid="24812" lane="2" />
                <ENTRY entrytime="NT" eventid="5686" heatid="24824" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Clara" gender="F" lastname="Schiller" nation="GER" license="420943" athleteid="24550">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.24" eventid="5712" heatid="24855" lane="3" />
                <ENTRY entrytime="00:01:12.92" eventid="5728" heatid="24871" lane="4" />
                <ENTRY entrytime="00:01:02.66" eventid="5744" heatid="24899" lane="2" />
                <ENTRY entrytime="00:00:50.00" eventid="7809" heatid="24919" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Elsa" gender="F" lastname="Schmaus" nation="GER" license="420936" athleteid="24555">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.15" eventid="5682" heatid="24817" lane="6" />
                <ENTRY entrytime="00:00:37.57" eventid="5698" heatid="24833" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5664" heatid="24808" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Cem Leon" gender="M" lastname="Schulze Döring" nation="GER" license="346286" athleteid="24559">
              <ENTRIES>
                <ENTRY entrytime="00:02:39.51" eventid="1177" heatid="24838" lane="2" />
                <ENTRY entrytime="00:00:42.26" eventid="5724" heatid="24870" lane="2" />
                <ENTRY entrytime="00:01:28.09" eventid="1165" heatid="24930" lane="2" />
                <ENTRY entrytime="00:03:06.56" eventid="5655" heatid="24947" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Finn Tolgar" gender="M" lastname="Schulze Döring" nation="GER" license="368690" athleteid="24783">
              <ENTRIES>
                <ENTRY entrytime="00:01:48.00" eventid="1141" heatid="24881" lane="6" />
                <ENTRY entrytime="00:01:58.00" eventid="7773" heatid="24908" lane="5" />
                <ENTRY entrytime="00:00:48.00" eventid="1117" heatid="24922" lane="3" />
                <ENTRY entrytime="00:01:32.94" eventid="1189" heatid="24936" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Nils Ömer" gender="M" lastname="Schulze Döring" nation="GER" license="393382" athleteid="24788">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.68" eventid="1053" heatid="24807" lane="3" />
                <ENTRY entrytime="00:00:21.63" eventid="5678" heatid="24814" lane="3" />
                <ENTRY entrytime="00:00:25.03" eventid="5694" heatid="24830" lane="3" />
                <ENTRY entrytime="00:00:00.30" eventid="7701" heatid="24834" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Julia" gender="F" lastname="Slonicz" nation="GER" license="430885" athleteid="23963">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.89" eventid="5664" heatid="24809" lane="2" />
                <ENTRY entrytime="00:00:39.55" eventid="5682" heatid="24817" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="5690" heatid="24828" lane="1" />
                <ENTRY entrytime="00:00:39.00" eventid="5698" heatid="24832" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-11-13" firstname="Tobias" gender="M" lastname="Steger" nation="GER" athleteid="24003">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.11" entrycourse="SCM" eventid="5702" heatid="24849" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.48" entrycourse="SCM" eventid="5724" heatid="24865" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.75" entrycourse="SCM" eventid="5740" heatid="24892" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-02-19" firstname="Nick" gender="M" lastname="Steinbinder" nation="GER" athleteid="24007">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.91" entrycourse="SCM" eventid="5702" heatid="24852" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.86" entrycourse="SCM" eventid="5740" heatid="24894" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="24935" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Roman" gender="M" lastname="Stroh" nation="GER" license="413758" athleteid="24793">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.87" eventid="5702" heatid="24849" lane="6" />
                <ENTRY entrytime="00:01:04.16" eventid="5724" heatid="24866" lane="1" />
                <ENTRY entrytime="00:01:02.44" eventid="5740" heatid="24890" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Amir" gender="M" lastname="Tawfik" nation="GER" license="420947" athleteid="24564">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="1053" heatid="24806" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5686" heatid="24825" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Annika" gender="F" lastname="Thummerer" nation="GER" license="393378" athleteid="24225">
              <ENTRIES>
                <ENTRY entrytime="00:04:00.00" eventid="1183" heatid="24840" lane="6" />
                <ENTRY entrytime="00:02:03.40" eventid="1135" heatid="24884" lane="3" />
                <ENTRY entrytime="00:02:15.28" eventid="7788" heatid="24911" lane="4" />
                <ENTRY entrytime="00:01:56.26" eventid="1195" heatid="24940" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jan" gender="M" lastname="Vilinski" nation="GER" athleteid="24567">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.00" eventid="5702" heatid="24848" lane="1" />
                <ENTRY entrytime="00:01:05.00" eventid="5724" heatid="24865" lane="3" />
                <ENTRY entrytime="00:01:02.00" eventid="5740" heatid="24891" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-04" firstname="Emily" gender="F" lastname="Wech" nation="GER" license="359178" athleteid="24011">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.07" entrycourse="SCM" eventid="1135" heatid="24886" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.74" entrycourse="SCM" eventid="7788" heatid="24914" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.71" entrycourse="SCM" eventid="1171" heatid="24931" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leander" gender="M" lastname="Wech" nation="GER" license="392571" athleteid="24571">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.85" eventid="5702" heatid="24848" lane="6" />
                <ENTRY entrytime="00:01:08.33" eventid="5724" heatid="24865" lane="1" />
                <ENTRY entrytime="00:01:02.39" eventid="5740" heatid="24890" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="7804" heatid="24917" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-10-19" firstname="Patrick" gender="M" lastname="Wech" nation="GER" license="392572" athleteid="24015">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.08" entrycourse="SCM" eventid="5724" heatid="24868" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.05" entrycourse="SCM" eventid="5740" heatid="24894" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.77" entrycourse="SCM" eventid="1117" heatid="24921" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Benjamin" gender="M" lastname="Welker" nation="GER" license="392569" athleteid="23968">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.56" eventid="5724" heatid="24866" lane="3" />
                <ENTRY entrytime="00:02:15.00" eventid="1141" heatid="24878" lane="4" />
                <ENTRY entrytime="00:00:25.00" eventid="7804" heatid="24918" lane="4" />
                <ENTRY entrytime="00:02:15.00" eventid="1189" heatid="24933" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Henri" gender="M" lastname="Wittl" nation="GER" athleteid="23973">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1053" heatid="24805" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="7691" heatid="24819" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="24825" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="F" lastname="Wolf" nation="GER" license="362947" athleteid="24576">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.15" eventid="1111" heatid="24863" lane="4" />
                <ENTRY entrytime="00:01:44.43" eventid="1135" heatid="24887" lane="3" />
                <ENTRY entrytime="00:01:32.82" eventid="7788" heatid="24916" lane="6" />
                <ENTRY entrytime="00:01:18.97" eventid="1195" heatid="24945" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Jan" gender="M" lastname="Zeidler" nation="GER" license="389378" athleteid="24797">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5702" heatid="24849" lane="5" />
                <ENTRY entrytime="NT" eventid="5724" heatid="24864" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="24891" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2015-01-01" firstname="Simon" gender="M" lastname="Zeidler" nation="GER" license="0" athleteid="24801">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.27" eventid="1053" heatid="24805" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5678" heatid="24813" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="24825" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-04-24" firstname="Arijalda" gender="F" lastname="Zukorlic" nation="GER" athleteid="24019">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="24853" lane="2" />
                <ENTRY entrytime="NT" eventid="5728" heatid="24871" lane="1" />
                <ENTRY entrytime="NT" eventid="5744" heatid="24898" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5085" nation="GER" region="02" clubid="24333" name="SG Bamberg">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="Elias" gender="M" lastname="Becker" nation="GER" license="429038" athleteid="24334">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="5702" heatid="24846" lane="4" />
                <ENTRY entrytime="00:01:20.00" eventid="5740" heatid="24889" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Katharina" gender="F" lastname="Dieter" nation="GER" license="0" athleteid="24337">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="24816" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="24821" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="24827" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Sanja" gender="F" lastname="Dietzel" nation="GER" license="0" athleteid="24341">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="24816" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="24822" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Mara" gender="F" lastname="Friedemann" nation="GER" license="434413" athleteid="24344">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.00" eventid="5712" heatid="24854" lane="6" />
                <ENTRY entrytime="00:01:30.00" eventid="5744" heatid="24898" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Leo" gender="M" lastname="Gebhard" nation="GER" license="425301" athleteid="24347">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.11" eventid="5702" heatid="24847" lane="1" />
                <ENTRY entrytime="00:01:10.00" eventid="5724" heatid="24865" lane="6" />
                <ENTRY entrytime="00:00:58.76" eventid="5740" heatid="24892" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Elisa" gender="F" lastname="Graf" nation="GER" license="0" athleteid="24351">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.94" eventid="5664" heatid="24808" lane="4" />
                <ENTRY entrytime="00:00:43.73" eventid="5682" heatid="24817" lane="1" />
                <ENTRY entrytime="00:00:55.00" eventid="7696" heatid="24822" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Emilia" gender="F" lastname="Graf" nation="GER" license="429036" athleteid="24355">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.00" eventid="5712" heatid="24854" lane="1" />
                <ENTRY entrytime="00:01:12.00" eventid="5728" heatid="24871" lane="3" />
                <ENTRY entrytime="00:01:06.00" eventid="5744" heatid="24899" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Moritz" gender="M" lastname="Hartmann" nation="GER" license="0" athleteid="24359">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.00" eventid="1053" heatid="24806" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5678" heatid="24813" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="7691" heatid="24819" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="24824" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Juna" gender="F" lastname="Heinze" nation="GER" license="0" athleteid="24364">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="24816" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Paula" gender="F" lastname="Heinze" nation="GER" license="395455" athleteid="24366">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.00" eventid="5712" heatid="24854" lane="3" />
                <ENTRY entrytime="00:01:09.00" eventid="5728" heatid="24872" lane="5" />
                <ENTRY entrytime="00:00:59.10" eventid="5744" heatid="24900" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Jannik" gender="M" lastname="Hünniger" nation="GER" license="409224" athleteid="24370">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.78" eventid="5702" heatid="24851" lane="2" />
                <ENTRY entrytime="00:00:47.54" eventid="5724" heatid="24869" lane="2" />
                <ENTRY entrytime="00:01:41.37" eventid="7773" heatid="24909" lane="1" />
                <ENTRY entrytime="00:01:46.00" eventid="1165" heatid="24929" lane="3" />
                <ENTRY entrytime="00:01:30.99" eventid="1189" heatid="24937" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lara" gender="F" lastname="Hünniger" nation="GER" license="425312" athleteid="24376">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.00" eventid="5712" heatid="24854" lane="5" />
                <ENTRY entrytime="00:00:59.20" eventid="5744" heatid="24900" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Timurs" gender="M" lastname="Iljins" nation="GER" license="409220" athleteid="24379">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="5702" heatid="24846" lane="3" />
                <ENTRY entrytime="00:00:58.88" eventid="5724" heatid="24866" lane="4" />
                <ENTRY entrytime="00:00:48.93" eventid="5740" heatid="24892" lane="3" />
                <ENTRY entrytime="00:02:15.00" eventid="7773" heatid="24907" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Eva" gender="F" lastname="Jakubaß" nation="GER" license="409223" athleteid="24384">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.80" eventid="5712" heatid="24855" lane="5" />
                <ENTRY entrytime="00:00:55.18" eventid="5728" heatid="24875" lane="1" />
                <ENTRY entrytime="00:00:48.65" eventid="5744" heatid="24902" lane="5" />
                <ENTRY entrytime="00:01:48.08" eventid="1195" heatid="24941" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Raphael" gender="M" lastname="Jakubaß" nation="GER" license="392827" athleteid="24389">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.99" eventid="5702" heatid="24849" lane="2" />
                <ENTRY entrytime="00:00:43.27" eventid="5740" heatid="24894" lane="4" />
                <ENTRY entrytime="00:01:50.00" eventid="7773" heatid="24908" lane="2" />
                <ENTRY entrytime="00:00:48.70" eventid="1117" heatid="24922" lane="4" />
                <ENTRY entrytime="00:01:39.77" eventid="1189" heatid="24936" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Sebastian" gender="M" lastname="Jakubaß" nation="GER" license="0" athleteid="24395">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5678" heatid="24812" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="7691" heatid="24819" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="24824" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Antonio" gender="M" lastname="La Corte" nation="GER" license="0" athleteid="24399">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5678" heatid="24812" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="24825" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Olivia" gender="F" lastname="Lang" nation="GER" license="425304" athleteid="24402">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5728" heatid="24872" lane="1" />
                <ENTRY entrytime="00:01:01.82" eventid="5744" heatid="24899" lane="3" />
                <ENTRY entrytime="00:00:36.00" eventid="7809" heatid="24920" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Samuel" gender="M" lastname="Lang" nation="GER" license="392828" athleteid="24406">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.00" eventid="1177" heatid="24837" lane="5" />
                <ENTRY entrytime="00:01:46.84" eventid="1103" heatid="24860" lane="4" />
                <ENTRY entrytime="00:00:37.28" eventid="5740" heatid="24896" lane="2" />
                <ENTRY entrytime="00:00:44.10" eventid="1117" heatid="24923" lane="5" />
                <ENTRY entrytime="00:01:25.60" eventid="1189" heatid="24937" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Eva" gender="F" lastname="Meister" nation="GER" license="409222" athleteid="24412">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.62" eventid="5712" heatid="24858" lane="6" />
                <ENTRY entrytime="00:01:02.76" eventid="5728" heatid="24873" lane="6" />
                <ENTRY entrytime="00:00:48.90" eventid="5744" heatid="24902" lane="6" />
                <ENTRY entrytime="00:02:07.00" eventid="7788" heatid="24912" lane="1" />
                <ENTRY entrytime="00:00:32.00" eventid="7809" heatid="24920" lane="1" />
                <ENTRY entrytime="00:01:55.00" eventid="1195" heatid="24940" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Jakob" gender="M" lastname="Meister" nation="GER" license="361866" athleteid="24419">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.00" eventid="5702" heatid="24852" lane="1" />
                <ENTRY entrytime="00:00:45.00" eventid="5724" heatid="24870" lane="1" />
                <ENTRY entrytime="00:00:38.00" eventid="5740" heatid="24896" lane="5" />
                <ENTRY entrytime="00:00:47.00" eventid="1117" heatid="24923" lane="6" />
                <ENTRY entrytime="00:01:39.00" eventid="1165" heatid="24930" lane="6" />
                <ENTRY entrytime="00:03:30.00" eventid="5655" heatid="24946" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Paul" gender="M" lastname="Nitsche" nation="GER" license="434412" athleteid="24426">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.00" eventid="5702" heatid="24846" lane="5" />
                <ENTRY entrytime="00:01:30.00" eventid="5740" heatid="24889" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Noa-Louis" gender="M" lastname="Panknin" nation="GER" license="429039" athleteid="24429">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5702" heatid="24847" lane="5" />
                <ENTRY entrytime="00:01:10.00" eventid="5740" heatid="24890" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Linda" gender="F" lastname="Schellenberger" nation="GER" license="0" athleteid="24432">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.00" eventid="5674" heatid="24811" lane="3" />
                <ENTRY entrytime="00:00:24.92" eventid="5682" heatid="24818" lane="3" />
                <ENTRY entrytime="00:00:29.10" eventid="7696" heatid="24823" lane="3" />
                <ENTRY entrytime="00:00:28.25" eventid="5698" heatid="24833" lane="3" />
                <ENTRY entrytime="00:00:36.00" eventid="7706" heatid="24835" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Marie" gender="F" lastname="Schellenberger" nation="GER" license="0" athleteid="24438">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.40" eventid="5664" heatid="24810" lane="4" />
                <ENTRY entrytime="00:00:33.06" eventid="5682" heatid="24818" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" heatid="24822" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="5690" heatid="24827" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lara" gender="F" lastname="Schindler" nation="GER" license="409221" athleteid="24443">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.26" eventid="5712" heatid="24857" lane="2" />
                <ENTRY entrytime="00:00:59.28" eventid="5728" heatid="24874" lane="4" />
                <ENTRY entrytime="00:00:52.03" eventid="5744" heatid="24901" lane="5" />
                <ENTRY entrytime="00:02:07.00" eventid="7788" heatid="24912" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Luisa" gender="F" lastname="Schindler" nation="GER" license="0" athleteid="24448">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5664" heatid="24808" lane="2" />
                <ENTRY entrytime="00:00:57.46" eventid="5682" heatid="24816" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="24822" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Paula" gender="F" lastname="Schuh" nation="GER" license="425299" athleteid="24452">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.11" eventid="5712" heatid="24855" lane="4" />
                <ENTRY entrytime="00:01:09.00" eventid="5728" heatid="24872" lane="2" />
                <ENTRY entrytime="00:00:56.49" eventid="5744" heatid="24900" lane="5" />
                <ENTRY entrytime="00:02:10.00" eventid="7788" heatid="24912" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Hanna" gender="F" lastname="Skamrahl" nation="GER" license="0" athleteid="24457">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5664" heatid="24808" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="24815" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="24827" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Antonia" gender="F" lastname="Struckmeier" nation="GER" license="0" athleteid="24461">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.36" eventid="5664" heatid="24809" lane="6" />
                <ENTRY entrytime="00:00:44.00" eventid="5674" heatid="24811" lane="4" />
                <ENTRY entrytime="00:00:32.20" eventid="5682" heatid="24818" lane="1" />
                <ENTRY entrytime="00:00:36.90" eventid="7696" heatid="24823" lane="4" />
                <ENTRY entrytime="00:00:41.34" eventid="5698" heatid="24832" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Troll" nation="GER" license="0" athleteid="24467">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5664" heatid="24808" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="24815" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="24822" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lilia" gender="F" lastname="Wagner" nation="GER" license="0" athleteid="24471">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="24816" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="24821" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="24827" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Laurin" gender="M" lastname="Willenberg" nation="GER" license="430362" athleteid="24475">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="5702" heatid="24847" lane="6" />
                <ENTRY entrytime="00:01:20.00" eventid="5740" heatid="24890" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Fiona" gender="F" lastname="Wystrach" nation="GER" license="0" athleteid="24478">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="24815" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="24821" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="24827" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5095" nation="GER" region="02" clubid="24581" name="SG Frankenhöhe">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="Laura" gender="F" lastname="Bauereiß" nation="GER" license="000000" athleteid="24582">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.00" eventid="5712" heatid="24857" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="24874" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5744" heatid="24901" lane="2" />
                <ENTRY entrytime="NT" eventid="7809" heatid="24919" lane="5" />
                <ENTRY entrytime="00:02:10.00" eventid="1195" heatid="24939" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Noah" gender="M" lastname="Binder" nation="GER" license="000000" athleteid="24588">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.00" eventid="5702" heatid="24851" lane="1" />
                <ENTRY entrytime="00:00:54.00" eventid="5724" heatid="24868" lane="5" />
                <ENTRY entrytime="00:00:39.00" eventid="5740" heatid="24895" lane="4" />
                <ENTRY entrytime="00:00:55.00" eventid="1117" heatid="24922" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Antonia" gender="F" lastname="Bößendorfer" nation="GER" license="364988" athleteid="24593">
              <ENTRIES>
                <ENTRY entrytime="00:03:01.27" eventid="1183" heatid="24844" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="1135" heatid="24886" lane="3" />
                <ENTRY entrytime="00:00:37.00" eventid="5744" heatid="24905" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="1123" heatid="24927" lane="1" />
                <ENTRY entrytime="00:01:25.00" eventid="1195" heatid="24944" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Emely" gender="F" lastname="Bößendörfer" nation="GER" license="364989" athleteid="24599">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.00" eventid="1183" heatid="24844" lane="4" />
                <ENTRY entrytime="00:01:40.00" eventid="1135" heatid="24888" lane="1" />
                <ENTRY entrytime="00:00:36.00" eventid="5744" heatid="24906" lane="5" />
                <ENTRY entrytime="00:00:44.00" eventid="1123" heatid="24928" lane="2" />
                <ENTRY entrytime="00:01:23.00" eventid="1195" heatid="24944" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Anne" gender="F" lastname="Frank" nation="GER" license="000000" athleteid="24605">
              <ENTRIES>
                <ENTRY entrytime="00:03:22.00" eventid="1183" heatid="24843" lane="2" />
                <ENTRY entrytime="00:01:49.00" eventid="1135" heatid="24887" lane="1" />
                <ENTRY entrytime="00:00:39.00" eventid="5744" heatid="24905" lane="5" />
                <ENTRY entrytime="00:00:55.00" eventid="1123" heatid="24926" lane="1" />
                <ENTRY entrytime="00:01:34.00" eventid="1195" heatid="24942" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lana" gender="F" lastname="Freisler" nation="GER" license="392397" athleteid="24611">
              <ENTRIES>
                <ENTRY entrytime="00:03:14.00" eventid="1183" heatid="24844" lane="6" />
                <ENTRY entrytime="00:01:45.00" eventid="1135" heatid="24887" lane="4" />
                <ENTRY entrytime="00:00:41.00" eventid="5744" heatid="24904" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="1123" heatid="24927" lane="5" />
                <ENTRY entrytime="00:01:32.00" eventid="1195" heatid="24943" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Jonah" gender="M" lastname="Henninger" nation="GER" license="379527" athleteid="24617">
              <ENTRIES>
                <ENTRY entrytime="00:02:25.00" eventid="1177" heatid="24838" lane="3" />
                <ENTRY entrytime="00:01:20.00" eventid="1103" heatid="24861" lane="3" />
                <ENTRY entrytime="00:00:29.00" eventid="5740" heatid="24897" lane="3" />
                <ENTRY entrytime="00:01:24.00" eventid="1165" heatid="24930" lane="4" />
                <ENTRY entrytime="00:01:05.00" eventid="1189" heatid="24938" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lea" gender="F" lastname="Herrmann" nation="GER" license="000000" athleteid="24623">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.00" eventid="5712" heatid="24857" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="24874" lane="5" />
                <ENTRY entrytime="00:00:49.00" eventid="5744" heatid="24901" lane="3" />
                <ENTRY entrytime="NT" eventid="7809" heatid="24919" lane="2" />
                <ENTRY entrytime="00:01:55.00" eventid="1195" heatid="24940" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Hanna" gender="F" lastname="Kachelrieß" nation="GER" license="392395" athleteid="24629">
              <ENTRIES>
                <ENTRY entrytime="00:03:25.00" eventid="1183" heatid="24843" lane="6" />
                <ENTRY entrytime="00:01:51.00" eventid="1135" heatid="24886" lane="4" />
                <ENTRY entrytime="00:00:39.00" eventid="5744" heatid="24905" lane="1" />
                <ENTRY entrytime="00:00:55.00" eventid="1123" heatid="24926" lane="6" />
                <ENTRY entrytime="00:01:31.00" eventid="1195" heatid="24943" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Julia" gender="F" lastname="KLaußecker" nation="GER" license="000000" athleteid="24635">
              <ENTRIES>
                <ENTRY entrytime="00:04:00.00" eventid="1183" heatid="24840" lane="1" />
                <ENTRY entrytime="00:01:55.00" eventid="1135" heatid="24886" lane="1" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="24901" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Sophia" gender="F" lastname="Kloha" nation="GER" license="000000" athleteid="24639">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.00" eventid="5712" heatid="24856" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="24873" lane="4" />
                <ENTRY entrytime="00:00:49.00" eventid="5744" heatid="24901" lane="4" />
                <ENTRY entrytime="00:01:55.00" eventid="1195" heatid="24941" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Eleni" gender="F" lastname="Martin" nation="GER" license="000000" athleteid="24644">
              <ENTRIES>
                <ENTRY entrytime="00:03:35.00" eventid="1183" heatid="24841" lane="3" />
                <ENTRY entrytime="00:01:55.00" eventid="1135" heatid="24886" lane="5" />
                <ENTRY entrytime="00:00:40.00" eventid="5744" heatid="24904" lane="3" />
                <ENTRY entrytime="00:01:38.00" eventid="1195" heatid="24942" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Eileen" gender="F" lastname="Möhring" nation="GER" license="000000" athleteid="24649">
              <ENTRIES>
                <ENTRY entrytime="00:02:58.00" eventid="1183" heatid="24845" lane="1" />
                <ENTRY entrytime="00:00:48.00" eventid="5728" heatid="24876" lane="4" />
                <ENTRY entrytime="00:00:36.00" eventid="5744" heatid="24906" lane="2" />
                <ENTRY entrytime="00:01:25.00" eventid="1195" heatid="24944" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Tilly" gender="F" lastname="Neumeyer" nation="GER" license="000000" athleteid="24654">
              <ENTRIES>
                <ENTRY entrytime="00:03:50.00" eventid="1183" heatid="24841" lane="6" />
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="24885" lane="6" />
                <ENTRY entrytime="00:00:45.00" eventid="5744" heatid="24903" lane="6" />
                <ENTRY entrytime="00:01:50.00" eventid="1195" heatid="24941" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Laurens" gender="M" lastname="Springer" nation="GER" license="000000" athleteid="24659">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.00" eventid="5702" heatid="24848" lane="5" />
                <ENTRY entrytime="00:01:08.00" eventid="5724" heatid="24865" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5740" heatid="24892" lane="4" />
                <ENTRY entrytime="00:01:55.00" eventid="1189" heatid="24934" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6621" nation="GER" region="02" clubid="24230" name="SG Rödental">
          <ATHLETES>
            <ATHLETE birthdate="2010-01-01" firstname="Esther" gender="F" lastname="Amberg" nation="GER" license="420966" athleteid="24231">
              <ENTRIES>
                <ENTRY entrytime="00:03:55.00" eventid="1183" heatid="24840" lane="2" />
                <ENTRY entrytime="00:00:55.62" eventid="5728" heatid="24875" lane="6" />
                <ENTRY entrytime="00:02:04.51" eventid="7788" heatid="24912" lane="3" />
                <ENTRY entrytime="00:00:32.00" eventid="7809" heatid="24920" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Theresa" gender="F" lastname="Dressel" nation="GER" license="0" athleteid="24236">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.00" eventid="5664" heatid="24810" lane="5" />
                <ENTRY entrytime="00:00:43.00" eventid="5682" heatid="24817" lane="5" />
                <ENTRY entrytime="00:00:39.00" eventid="5690" heatid="24828" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="24831" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Hannes" gender="M" lastname="Endruweit" nation="GER" license="0" athleteid="24241">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="1053" heatid="24806" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="5678" heatid="24814" lane="6" />
                <ENTRY entrytime="00:00:35.00" eventid="7691" heatid="24820" lane="3" />
                <ENTRY entrytime="00:00:55.00" eventid="7701" heatid="24834" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Jannik" gender="M" lastname="Endruweit" nation="GER" license="380996" athleteid="24246">
              <ENTRIES>
                <ENTRY entrytime="00:02:48.61" eventid="1177" heatid="24838" lane="5" />
                <ENTRY entrytime="00:01:29.55" eventid="1103" heatid="24861" lane="2" />
                <ENTRY entrytime="00:01:27.58" eventid="7773" heatid="24910" lane="5" />
                <ENTRY entrytime="00:00:18.00" eventid="7804" heatid="24918" lane="3" />
                <ENTRY entrytime="00:01:15.20" eventid="1189" heatid="24938" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Emely" gender="F" lastname="Gräser" nation="GER" license="367553" athleteid="24252">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.42" eventid="5728" heatid="24877" lane="3" />
                <ENTRY entrytime="00:00:34.05" eventid="5744" heatid="24906" lane="3" />
                <ENTRY entrytime="00:01:28.86" eventid="7788" heatid="24916" lane="4" />
                <ENTRY entrytime="00:01:23.08" eventid="1171" heatid="24932" lane="3" />
                <ENTRY entrytime="00:01:14.45" eventid="1195" heatid="24945" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Till" gender="M" lastname="Gräser" nation="GER" license="404231" athleteid="24258">
              <ENTRIES>
                <ENTRY entrytime="00:03:36.42" eventid="1177" heatid="24836" lane="4" />
                <ENTRY entrytime="00:00:48.88" eventid="5724" heatid="24869" lane="5" />
                <ENTRY entrytime="00:00:38.51" eventid="5740" heatid="24896" lane="6" />
                <ENTRY entrytime="00:00:30.00" eventid="7804" heatid="24917" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Anne-Lotte" gender="F" lastname="Hofbauer" nation="GER" license="417943" athleteid="24263">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.70" eventid="5712" heatid="24856" lane="1" />
                <ENTRY entrytime="00:02:19.64" eventid="1135" heatid="24882" lane="3" />
                <ENTRY entrytime="00:00:47.02" eventid="5744" heatid="24902" lane="2" />
                <ENTRY entrytime="00:02:10.00" eventid="1171" heatid="24931" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lennart" gender="M" lastname="Hofbauer" nation="GER" license="364856" athleteid="24268">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.44" eventid="5702" heatid="24852" lane="4" />
                <ENTRY entrytime="00:00:46.66" eventid="5724" heatid="24869" lane="3" />
                <ENTRY entrytime="00:00:33.97" eventid="5740" heatid="24897" lane="1" />
                <ENTRY entrytime="00:01:33.00" eventid="7773" heatid="24910" lane="6" />
                <ENTRY entrytime="00:01:14.96" eventid="1189" heatid="24938" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Jonathan" gender="M" lastname="Kohles" nation="GER" license="373339" athleteid="24274">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.83" eventid="1103" heatid="24861" lane="5" />
                <ENTRY entrytime="00:01:23.99" eventid="1141" heatid="24881" lane="3" />
                <ENTRY entrytime="00:01:22.00" eventid="7773" heatid="24910" lane="4" />
                <ENTRY entrytime="00:00:37.00" eventid="1117" heatid="24923" lane="3" />
                <ENTRY entrytime="00:01:13.89" eventid="1189" heatid="24938" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Sophia" gender="F" lastname="Lamik" nation="GER" license="0" athleteid="24280">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.00" eventid="5664" heatid="24809" lane="5" />
                <ENTRY entrytime="00:00:42.00" eventid="7696" heatid="24823" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="24832" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="7706" heatid="24835" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Arne" gender="M" lastname="Mesch" nation="GER" license="361790" athleteid="24285">
              <ENTRIES>
                <ENTRY entrytime="00:02:33.29" eventid="1177" heatid="24838" lane="4" />
                <ENTRY entrytime="00:00:37.81" eventid="5724" heatid="24870" lane="4" />
                <ENTRY entrytime="00:01:19.61" eventid="7773" heatid="24910" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="1117" heatid="24923" lane="4" />
                <ENTRY entrytime="00:01:08.15" eventid="1189" heatid="24938" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Tobais Damian" gender="M" lastname="Schiebert" nation="GER" license="429408" athleteid="24291">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5702" heatid="24847" lane="2" />
                <ENTRY entrytime="00:01:10.00" eventid="5724" heatid="24864" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="24891" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Manuel" gender="M" lastname="Staffel" nation="GER" license="364847" athleteid="24295">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.41" eventid="1177" heatid="24838" lane="6" />
                <ENTRY entrytime="00:00:35.54" eventid="5740" heatid="24896" lane="3" />
                <ENTRY entrytime="00:01:38.64" eventid="7773" heatid="24909" lane="5" />
                <ENTRY entrytime="00:01:38.02" eventid="1165" heatid="24930" lane="1" />
                <ENTRY entrytime="00:01:17.76" eventid="1189" heatid="24937" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lea" gender="F" lastname="Tarrach" nation="GER" license="373337" athleteid="24301">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.25" eventid="5712" heatid="24859" lane="3" />
                <ENTRY entrytime="00:01:34.79" eventid="1135" heatid="24888" lane="3" />
                <ENTRY entrytime="00:00:36.21" eventid="5744" heatid="24906" lane="1" />
                <ENTRY entrytime="00:01:38.00" eventid="7788" heatid="24915" lane="2" />
                <ENTRY entrytime="00:01:21.11" eventid="1195" heatid="24944" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lina" gender="F" lastname="Tarrach" nation="GER" license="417942" athleteid="24307">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.39" eventid="5712" heatid="24857" lane="5" />
                <ENTRY entrytime="00:01:02.40" eventid="5728" heatid="24873" lane="1" />
                <ENTRY entrytime="00:02:07.72" eventid="1135" heatid="24884" lane="6" />
                <ENTRY entrytime="00:02:05.00" eventid="1195" heatid="24939" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Johanna" gender="F" lastname="Thiem" nation="GER" license="404230" athleteid="24312">
              <ENTRIES>
                <ENTRY entrytime="00:03:33.93" eventid="1183" heatid="24842" lane="6" />
                <ENTRY entrytime="00:01:59.86" eventid="7788" heatid="24913" lane="2" />
                <ENTRY entrytime="00:00:50.56" eventid="1123" heatid="24926" lane="3" />
                <ENTRY entrytime="00:01:48.13" eventid="1195" heatid="24941" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Vanessa" gender="F" lastname="Thiem" nation="GER" license="404232" athleteid="24317">
              <ENTRIES>
                <ENTRY entrytime="00:02:57.28" eventid="1183" heatid="24845" lane="5" />
                <ENTRY entrytime="00:00:35.95" eventid="5744" heatid="24906" lane="4" />
                <ENTRY entrytime="00:01:34.05" eventid="7788" heatid="24915" lane="3" />
                <ENTRY entrytime="00:00:42.81" eventid="1123" heatid="24928" lane="3" />
                <ENTRY entrytime="00:01:19.53" eventid="1195" heatid="24945" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Alina" gender="F" lastname="Zeder" nation="GER" license="0" athleteid="24323">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.00" eventid="5664" heatid="24809" lane="4" />
                <ENTRY entrytime="00:00:39.00" eventid="7696" heatid="24823" lane="2" />
                <ENTRY entrytime="00:00:37.00" eventid="5690" heatid="24828" lane="2" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="24832" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Bastian" gender="M" lastname="Zetzmann" nation="GER" license="392527" athleteid="24328">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.55" eventid="5702" heatid="24850" lane="2" />
                <ENTRY entrytime="00:02:00.73" eventid="1141" heatid="24880" lane="1" />
                <ENTRY entrytime="00:02:05.00" eventid="7773" heatid="24907" lane="3" />
                <ENTRY entrytime="00:01:48.00" eventid="1189" heatid="24935" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4502" nation="GER" region="02" clubid="24023" name="TSV Zirndorf">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Jana" gender="F" lastname="Ammon" nation="GER" license="398728" athleteid="24024">
              <ENTRIES>
                <ENTRY entrytime="00:03:00.00" eventid="1183" heatid="24845" lane="6" />
                <ENTRY entrytime="00:01:40.00" eventid="1111" heatid="24863" lane="2" />
                <ENTRY entrytime="00:00:41.63" eventid="5744" heatid="24903" lane="4" />
                <ENTRY entrytime="00:01:46.09" eventid="1171" heatid="24932" lane="5" />
                <ENTRY entrytime="00:01:27.68" eventid="1195" heatid="24944" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Marco" gender="M" lastname="Ammon" nation="GER" license="398727" athleteid="24030">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.00" eventid="1177" heatid="24838" lane="1" />
                <ENTRY entrytime="00:01:48.15" eventid="1141" heatid="24880" lane="3" />
                <ENTRY entrytime="00:01:38.56" eventid="7773" heatid="24909" lane="2" />
                <ENTRY entrytime="00:00:46.85" eventid="1117" heatid="24923" lane="1" />
                <ENTRY entrytime="00:02:50.00" eventid="5655" heatid="24947" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Alissa" gender="F" lastname="Bader" nation="GER" license="428030" athleteid="24036">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.00" eventid="1183" heatid="24844" lane="1" />
                <ENTRY entrytime="00:00:50.28" eventid="5712" heatid="24859" lane="6" />
                <ENTRY entrytime="00:01:56.25" eventid="1135" heatid="24886" lane="6" />
                <ENTRY entrytime="00:00:40.06" eventid="5744" heatid="24904" lane="4" />
                <ENTRY entrytime="00:01:36.53" eventid="1195" heatid="24942" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Mia" gender="F" lastname="Großhauser" nation="GER" license="420483" athleteid="24042">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.00" eventid="1183" heatid="24844" lane="5" />
                <ENTRY entrytime="00:01:59.09" eventid="1135" heatid="24885" lane="1" />
                <ENTRY entrytime="00:01:53.94" eventid="7788" heatid="24913" lane="3" />
                <ENTRY entrytime="00:00:25.12" eventid="7809" heatid="24920" lane="3" />
                <ENTRY entrytime="00:01:35.78" eventid="1195" heatid="24942" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Josefine" gender="F" lastname="Mendler" nation="GER" license="420484" athleteid="24048">
              <ENTRIES>
                <ENTRY entrytime="00:03:40.00" eventid="1183" heatid="24841" lane="5" />
                <ENTRY entrytime="00:01:08.35" eventid="5728" heatid="24872" lane="4" />
                <ENTRY entrytime="00:02:08.52" eventid="1135" heatid="24883" lane="3" />
                <ENTRY entrytime="00:02:05.00" eventid="7788" heatid="24912" lane="4" />
                <ENTRY entrytime="00:02:02.26" eventid="1195" heatid="24940" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Simona" gender="F" lastname="Paschold" nation="GER" license="398731" athleteid="24054">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.74" eventid="1183" heatid="24845" lane="4" />
                <ENTRY entrytime="00:00:45.09" eventid="5728" heatid="24877" lane="1" />
                <ENTRY entrytime="00:01:37.69" eventid="1135" heatid="24888" lane="4" />
                <ENTRY entrytime="00:01:30.12" eventid="7788" heatid="24916" lane="5" />
                <ENTRY entrytime="00:00:45.56" eventid="1123" heatid="24928" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Tim Simon" gender="M" lastname="Paschold" nation="GER" license="428031" athleteid="24060">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.50" eventid="5702" heatid="24848" lane="4" />
                <ENTRY entrytime="00:01:05.93" eventid="5724" heatid="24865" lane="2" />
                <ENTRY entrytime="00:02:14.09" eventid="1141" heatid="24878" lane="3" />
                <ENTRY entrytime="00:00:48.87" eventid="5740" heatid="24893" lane="6" />
                <ENTRY entrytime="00:02:00.56" eventid="1189" heatid="24934" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
