<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SG Fürth" version="11.61084">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Nürnberg" name="Bayerische Kurzbahnmeisterschaften 2019" course="SCM" deadline="2016-10-26" hostclub="SG Mittelfranken" organizer="Bayerischer Schwimmverband e.V." organizer.url="http://www.bayerischer-schwimmverband.de/schwimmen" reservecount="4" startmethod="1" timing="AUTOMATIC" nation="GER">
      <AGEDATE value="2016-11-06" type="YEAR" />
      <POOL name="90471 Nürnberg, Hallenbad Langwasser, Breslauer Str. 251, Eingang Gleiwitzer Straße" lanemin="1" lanemax="6" />
      <FACILITY city="Nürnberg" name="90471 Nürnberg, Hallenbad Langwasser, Breslauer Str. 251, Eingang Gleiwitzer Straße" nation="GER" />
      <POINTTABLE pointtableid="3009" name="FINA Point Scoring" version="2016" />
      <CONTACT city="Fürth" email="meldungen@sgfuerth.de" name="Matthias Fuchs" phone="09118101172" street="Lavendelweg 47" zip="90768" />
      <QUALIFY from="2016-01-01" until="2016-10-28" />
      <SESSIONS>
        <SESSION date="2016-11-05" daytime="10:00" number="1" officialmeeting="09:30" teamleadermeeting="09:30" warmupfrom="08:30" warmupuntil="09:50">
          <EVENTS>
            <EVENT eventid="1841" daytime="14:05" gender="F" number="15" order="26" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4779" daytime="14:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4780" daytime="14:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4781" daytime="14:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4782" daytime="14:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4783" daytime="14:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4784" daytime="14:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1763" daytime="10:50" gender="M" number="4" order="7" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4696" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4697" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4698" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4699" daytime="10:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4700" daytime="10:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4701" daytime="10:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4702" daytime="11:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4703" daytime="11:00" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1813" daytime="12:45" gender="F" number="11" order="19" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4745" daytime="12:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4746" daytime="12:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4747" daytime="12:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1792" daytime="11:50" gender="M" number="8" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4726" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4727" daytime="12:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1827" daytime="13:15" gender="F" number="13" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4758" daytime="13:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4759" daytime="13:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4760" daytime="13:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4761" daytime="13:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4762" daytime="13:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4763" daytime="13:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4764" daytime="13:50" number="7" order="7" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1820" daytime="12:55" gender="M" number="12" order="20" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4749" daytime="12:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4750" daytime="13:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4751" daytime="13:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4752" daytime="13:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4753" daytime="13:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4754" daytime="13:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4755" daytime="13:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4756" daytime="13:15" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1756" daytime="10:40" gender="F" number="3" order="5" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4687" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4688" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4689" daytime="10:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4690" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4691" daytime="10:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4692" daytime="10:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4693" daytime="10:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4694" daytime="10:45" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1785" daytime="11:40" gender="F" number="7" order="13" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4718" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4719" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4720" daytime="11:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4721" daytime="11:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4722" daytime="11:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4723" daytime="11:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4724" daytime="11:45" number="7" order="7" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1749" daytime="10:20" gender="M" number="2" order="3" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4676" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4677" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4678" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4679" daytime="10:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4680" daytime="10:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4681" daytime="10:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4682" daytime="10:30" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4683" daytime="10:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4684" daytime="10:35" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4685" daytime="10:40" number="10" order="10" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1806" daytime="12:40" gender="M" number="10" order="18" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4738" daytime="12:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4739" daytime="12:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4740" daytime="12:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4741" daytime="12:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4742" daytime="12:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4743" daytime="12:45" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1778" daytime="11:25" gender="M" number="6" order="11" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4709" daytime="11:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4710" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4711" daytime="11:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4712" daytime="11:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4713" daytime="11:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4714" daytime="11:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4715" daytime="11:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4716" daytime="11:35" number="8" order="8" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5369" gender="M" number="6" order="30" round="SOP" preveventid="1778">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="5378" agegroupid="5375" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1059" daytime="10:00" gender="F" number="1" order="1" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4662" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4663" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4664" daytime="10:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4665" daytime="10:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4666" daytime="10:05" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4667" daytime="10:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4668" daytime="10:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4669" daytime="10:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4670" daytime="10:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4671" daytime="10:10" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4672" daytime="10:15" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4673" daytime="10:15" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4674" daytime="10:15" number="13" order="13" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5443" gender="M" number="14" order="31" round="SOP" preveventid="1834">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="5452" agegroupid="5449" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1848" daytime="14:25" gender="M" number="16" order="27" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4786" daytime="14:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4787" daytime="14:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4788" daytime="14:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4789" daytime="14:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4790" daytime="14:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4791" daytime="14:35" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1771" daytime="11:00" gender="F" number="5" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4705" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4706" daytime="11:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4707" daytime="11:15" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4708" daytime="11:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1855" daytime="14:40" gender="F" number="17" order="28" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4793" daytime="14:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4794" daytime="14:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4795" daytime="14:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4796" daytime="14:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4797" daytime="14:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4798" daytime="14:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4799" daytime="14:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4800" daytime="14:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4801" daytime="14:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4961" daytime="14:45" number="10" order="10" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1799" daytime="12:25" gender="F" number="9" order="16" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4728" daytime="12:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4729" daytime="12:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4730" daytime="12:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4731" daytime="12:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4732" daytime="12:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4733" daytime="12:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4734" daytime="12:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4735" daytime="12:35" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4736" daytime="12:35" number="9" order="9" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1834" daytime="13:55" gender="M" number="14" order="24" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4765" daytime="13:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4766" daytime="13:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4767" daytime="13:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4768" daytime="13:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4769" daytime="13:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4770" daytime="13:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4771" daytime="13:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4772" daytime="14:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4773" daytime="14:00" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4774" daytime="14:00" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4775" daytime="14:00" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4776" daytime="14:00" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4777" daytime="14:00" number="13" order="13" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-11-05" daytime="16:45" endtime="19:39" number="2">
          <EVENTS>
            <EVENT eventid="1919" gender="F" number="9" order="25" round="FIN" preveventid="1799">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="5404" agegroupid="1920" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4737" agegroupid="1920" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1898" gender="M" number="6" order="18" round="FIN" preveventid="1778">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="5465" agegroupid="1899" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4717" agegroupid="1899" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1905" gender="F" number="18" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4803" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4804" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1863" gender="F" number="1" order="3" round="FIN" preveventid="1059">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="5317" agegroupid="1864" final="B" number="1" order="1" status="INOFFICIAL" />
                <HEAT heatid="4675" agegroupid="1864" final="A" number="2" order="2" status="INOFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1926" gender="M" number="12" order="27" round="FIN" preveventid="1820">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="5442" agegroupid="1927" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4757" agegroupid="1927" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1954" gender="F" number="15" order="33" round="FIN" preveventid="1841">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="5491" agegroupid="1955" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4785" agegroupid="1955" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1884" gender="M" number="4" order="13" round="FIN" preveventid="1763">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="5368" agegroupid="1885" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4704" agegroupid="1885" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2062" gender="F" number="20" order="41" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="2000" />
              <HEATS>
                <HEAT heatid="4807" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1870" gender="M" number="2" order="6" round="FIN" preveventid="1749">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="5342" agegroupid="1871" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4686" agegroupid="1871" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1891" gender="F" number="7" order="15" round="FIN" preveventid="1785">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="5391" agegroupid="1892" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4725" agegroupid="1892" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1912" gender="M" number="10" order="23" round="FIN" preveventid="1806">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="5417" agegroupid="1913" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4744" agegroupid="1913" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1947" gender="M" number="14" order="31" round="FIN" preveventid="1834">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="5478" agegroupid="1948" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4778" agegroupid="1948" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1961" gender="M" number="16" order="35" round="FIN" preveventid="1848">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="5504" agegroupid="1962" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4792" agegroupid="1962" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1877" gender="F" number="3" order="10" round="FIN" preveventid="1756">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="5355" agegroupid="1878" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4695" agegroupid="1878" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2048" gender="M" number="19" order="40" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="2000" />
              <HEATS>
                <HEAT heatid="4805" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4806" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1933" gender="F" number="11" order="29" round="FIN" preveventid="1813">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="5429" agegroupid="1934" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4748" agegroupid="1934" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1940" gender="F" number="17" order="37" round="FIN" preveventid="1855">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="5517" agegroupid="1941" final="B" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4802" agegroupid="1941" final="A" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-11-06" daytime="09:30" number="3" officialmeeting="09:00" teamleadermeeting="09:00" warmupfrom="07:45" warmupuntil="09:15">
          <EVENTS>
            <EVENT eventid="1999" daytime="10:35" gender="M" number="25" order="32" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4859" daytime="10:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4860" daytime="10:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4861" daytime="10:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4862" daytime="10:50" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1971" daytime="09:30" gender="M" number="21" order="23" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4813" daytime="09:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4814" daytime="09:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4815" daytime="09:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4816" daytime="09:35" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4817" daytime="09:35" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4818" daytime="09:35" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4819" daytime="09:35" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4820" daytime="09:40" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4821" daytime="09:40" number="9" order="9" status="SEEDED" />
                <HEAT heatid="4822" daytime="09:40" number="10" order="10" status="SEEDED" />
                <HEAT heatid="4823" daytime="09:40" number="11" order="11" status="SEEDED" />
                <HEAT heatid="4824" daytime="09:45" number="12" order="12" status="SEEDED" />
                <HEAT heatid="4825" daytime="09:45" number="13" order="13" status="SEEDED" />
                <HEAT heatid="4826" daytime="09:45" number="14" order="14" status="SEEDED" />
                <HEAT heatid="4827" daytime="09:45" number="15" order="15" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2096" daytime="13:30" gender="F" number="36" order="49" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4932" daytime="13:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4933" daytime="13:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4934" daytime="13:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4935" daytime="13:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4936" daytime="13:40" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4937" daytime="13:45" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1985" daytime="10:15" gender="M" number="23" order="28" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4840" daytime="10:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4841" daytime="10:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4842" daytime="10:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4843" daytime="10:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4844" daytime="10:20" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4845" daytime="10:20" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4846" daytime="10:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4847" daytime="10:20" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4848" daytime="10:20" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2027" daytime="11:35" gender="M" number="29" order="39" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4877" daytime="11:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4878" daytime="11:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4879" daytime="11:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4880" daytime="11:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4881" daytime="11:40" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2013" daytime="11:05" gender="M" number="27" order="36" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4869" daytime="11:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4870" daytime="11:10" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4871" daytime="11:10" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4872" daytime="11:10" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4873" daytime="11:10" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1978" daytime="09:50" gender="F" number="22" order="26" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4829" daytime="09:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4830" daytime="09:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4831" daytime="09:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4832" daytime="09:55" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4833" daytime="10:00" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4834" daytime="10:00" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4835" daytime="10:05" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4836" daytime="10:05" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4837" daytime="10:10" number="9" order="9" status="SEEDED" />
                <HEAT heatid="4838" daytime="10:10" number="10" order="10" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1992" daytime="10:20" gender="F" number="24" order="30" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4850" daytime="10:20" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4851" daytime="10:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4852" daytime="10:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4853" daytime="10:25" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4854" daytime="10:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4855" daytime="10:30" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4856" daytime="10:30" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4857" daytime="10:35" number="8" order="8" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2055" daytime="12:00" gender="F" number="32" order="43" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4896" daytime="12:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4897" daytime="12:05" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4898" daytime="12:10" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4899" daytime="12:10" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4900" daytime="12:15" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4901" daytime="12:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4902" daytime="12:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4903" daytime="12:20" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4904" daytime="12:25" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2075" daytime="12:30" gender="M" number="33" order="44" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4906" daytime="12:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4907" daytime="12:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4908" daytime="12:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4909" daytime="12:45" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4910" daytime="12:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4911" daytime="12:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4912" daytime="12:55" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2034" daytime="11:45" gender="F" number="30" order="41" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4883" daytime="11:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4884" daytime="11:45" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4885" daytime="11:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4886" daytime="11:45" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4887" daytime="11:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4888" daytime="11:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4889" daytime="11:50" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2103" daytime="13:45" gender="M" number="37" order="50" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4939" daytime="13:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4940" daytime="13:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4941" daytime="13:50" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4942" daytime="13:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4943" daytime="13:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4944" daytime="13:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4945" daytime="13:50" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4946" daytime="13:50" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4947" daytime="13:55" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2006" daytime="10:55" gender="F" number="26" order="34" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4863" daytime="10:55" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4864" daytime="11:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4865" daytime="11:00" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4866" daytime="11:00" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4867" daytime="11:05" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2041" daytime="11:50" gender="M" number="31" order="42" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4891" daytime="11:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4892" daytime="11:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4893" daytime="11:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4894" daytime="12:00" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2082" daytime="13:00" gender="F" number="34" order="46" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4913" daytime="13:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4914" daytime="13:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4915" daytime="13:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4916" daytime="13:05" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4917" daytime="13:05" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4918" daytime="13:05" number="6" order="6" status="SEEDED" />
                <HEAT heatid="4919" daytime="13:05" number="7" order="7" status="SEEDED" />
                <HEAT heatid="4920" daytime="13:05" number="8" order="8" status="SEEDED" />
                <HEAT heatid="4921" daytime="13:05" number="9" order="9" status="SEEDED" />
                <HEAT heatid="4922" daytime="13:10" number="10" order="10" status="SEEDED" />
                <HEAT heatid="4923" daytime="13:10" number="11" order="11" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2089" daytime="13:10" gender="M" number="35" order="48" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4925" daytime="13:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4926" daytime="13:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="4927" daytime="13:20" number="3" order="3" status="SEEDED" />
                <HEAT heatid="4928" daytime="13:20" number="4" order="4" status="SEEDED" />
                <HEAT heatid="4929" daytime="13:25" number="5" order="5" status="SEEDED" />
                <HEAT heatid="4930" daytime="13:25" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2020" daytime="11:15" gender="F" number="28" order="37" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4875" daytime="11:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4876" daytime="11:25" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2016-11-06" daytime="16:00" number="4">
          <EVENTS>
            <EVENT eventid="2154" gender="F" number="26" order="52" round="FIN" preveventid="2006">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="4868" agegroupid="2155" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2210" gender="M" number="35" order="70" round="FIN" preveventid="2089">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="4931" agegroupid="2211" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2168" gender="M" number="38" order="55" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="1000" />
              <HEATS>
                <HEAT heatid="4808" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4809" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2189" gender="M" number="31" order="66" round="FIN" preveventid="2041">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="4895" agegroupid="2190" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2182" gender="F" number="30" order="57" round="FIN" preveventid="2034">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="4890" agegroupid="2183" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2126" gender="M" number="21" order="41" round="FIN" preveventid="1971">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="4828" agegroupid="2127" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2147" gender="F" number="24" order="48" round="FIN" preveventid="1992">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="4858" agegroupid="2148" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2224" gender="F" number="39" order="77" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE value="2000" />
              <HEATS>
                <HEAT heatid="4810" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2133" gender="F" number="22" order="43" round="FIN" preveventid="1978">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="4839" agegroupid="2134" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2112" gender="M" number="37" order="74" round="FIN" preveventid="2103">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="4948" agegroupid="2113" final="A" number="1" order="1" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2175" gender="M" number="29" order="60" round="FIN" preveventid="2027">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="4882" agegroupid="2176" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2232" gender="M" number="40" order="78" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE value="2000" />
              <HEATS>
                <HEAT heatid="4811" number="1" order="1" status="SEEDED" />
                <HEAT heatid="4812" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="2070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2140" gender="M" number="23" order="46" round="FIN" preveventid="1985">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="4849" agegroupid="2141" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2203" gender="F" number="34" order="68" round="FIN" preveventid="2082">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="4924" agegroupid="2204" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2196" gender="F" number="32" order="64" round="FIN" preveventid="2055">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="4905" agegroupid="2197" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2217" gender="F" number="36" order="72" round="FIN" preveventid="2096">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="4938" agegroupid="2218" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1064" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2161" gender="M" number="27" order="50" round="FIN" preveventid="2013">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="4874" agegroupid="2162" final="A" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1066" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1078" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1070" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="4167" nation="GER" region="02" clubid="2398" name="1.SC Schweinfurt">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Daniel" gender="M" lastname="Heidbeck" nation="GER" license="379928" athleteid="2399">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.10" eventid="1763" heatid="4696" lane="4" />
                <ENTRY entrytime="00:00:34.57" eventid="1985" heatid="4841" lane="1" />
                <ENTRY entrytime="00:02:41.81" eventid="2089" heatid="4925" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Simon" gender="M" lastname="Vollert" nation="GER" license="331888" athleteid="2403">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.34" eventid="1834" heatid="4765" lane="3" />
                <ENTRY entrytime="00:00:34.74" eventid="1985" heatid="4840" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4175" nation="GER" region="02" clubid="2525" name="ASV 1860 Neumarkt">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Anika" gender="F" lastname="Jacksteit" nation="GER" license="266125" athleteid="2526">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.58" eventid="1059" heatid="4665" lane="4" />
                <ENTRY entrytime="00:01:13.24" eventid="1785" heatid="4718" lane="4" />
                <ENTRY entrytime="00:01:13.23" eventid="1799" heatid="4730" lane="5" />
                <ENTRY entrytime="00:00:33.63" eventid="2034" heatid="4885" lane="1" />
                <ENTRY entrytime="00:00:29.02" eventid="2082" heatid="4916" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4168" nation="GER" region="02" clubid="2759" name="ASV Cham">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Lena" gender="F" lastname="Braun" nation="GER" license="294440" athleteid="2760">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.92" eventid="1059" heatid="4670" lane="1" />
                <ENTRY entrytime="00:00:34.84" eventid="1756" heatid="4694" lane="6" />
                <ENTRY entrytime="00:01:12.36" eventid="1799" heatid="4732" lane="5" />
                <ENTRY entrytime="00:01:18.92" eventid="1992" heatid="4852" lane="3" />
                <ENTRY entrytime="00:00:27.35" eventid="2082" heatid="4921" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Alexandra" gender="F" lastname="Wagner" nation="GER" license="320557" athleteid="2766">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.10" eventid="1756" heatid="4688" lane="3" />
                <ENTRY entrytime="00:01:14.12" eventid="1799" heatid="4730" lane="6" />
                <ENTRY entrytime="00:00:32.15" eventid="1855" heatid="4793" lane="4" />
                <ENTRY entrytime="00:00:29.53" eventid="2082" heatid="4915" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4169" nation="GER" region="02" clubid="4644" name="ATS Kulmbach">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Franz" gender="M" lastname="Prell" nation="GER" license="297312" athleteid="4645">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.83" eventid="1749" heatid="4677" lane="1" />
                <ENTRY entrytime="00:04:40.20" eventid="2075" heatid="4906" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4224" nation="GER" region="02" clubid="3447" name="Delphin 77 Herzogenaurach">
          <ATHLETES>
            <ATHLETE birthdate="1992-01-01" firstname="Christian" gender="M" lastname="Ziebuhr" nation="GER" license="139641" athleteid="3448">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.50" eventid="1763" heatid="4700" lane="1" />
                <ENTRY entrytime="00:00:25.65" eventid="1834" heatid="4771" lane="5" />
                <ENTRY entrytime="00:00:31.35" eventid="1985" heatid="4845" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4233" nation="GER" region="02" clubid="3238" name="DJK Sportbund München">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Stefanie" gender="F" lastname="Ohneiser" nation="GER" license="316235" athleteid="3239">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.50" eventid="1059" heatid="4663" lane="4" />
                <ENTRY entrytime="00:01:15.00" eventid="1799" heatid="4728" lane="3" />
                <ENTRY entrytime="00:04:57.50" eventid="1827" heatid="4758" lane="2" />
                <ENTRY entrytime="00:00:31.00" eventid="1855" heatid="4797" lane="4" />
                <ENTRY entrytime="00:02:18.50" eventid="1978" heatid="4831" lane="4" />
                <ENTRY entrytime="00:02:38.50" eventid="2055" heatid="4898" lane="6" />
                <ENTRY entrytime="00:00:29.50" eventid="2082" heatid="4915" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4300" nation="GER" region="02" clubid="2665" name="SB Bayern 07">
          <ATHLETES>
            <ATHLETE birthdate="1995-01-01" firstname="Tim" gender="M" lastname="Grasser" nation="GER" license="150609" athleteid="2666">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.90" eventid="1834" heatid="4770" lane="4" />
                <ENTRY entrytime="00:00:56.19" eventid="1971" heatid="4821" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Teresa" gender="F" lastname="Kraus" nation="GER" license="183593" athleteid="2669">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.29" eventid="1799" heatid="4732" lane="4" />
                <ENTRY entrytime="00:00:29.68" eventid="1855" heatid="4961" lane="1" />
                <ENTRY entrytime="00:01:08.50" eventid="2006" heatid="4864" lane="3" />
                <ENTRY entrytime="00:00:29.00" eventid="2082" heatid="4917" lane="6" />
                <ENTRY entrytime="00:01:10.47" eventid="1919" heatid="5404" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.42" eventid="1940" heatid="5517" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4290" nation="GER" region="02" clubid="2598" name="SC 53 Landshut">
          <ATHLETES>
            <ATHLETE birthdate="1993-01-01" firstname="Verena" gender="F" lastname="Dormehl" nation="GER" license="154254" athleteid="2599">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.45" eventid="1756" heatid="4691" lane="4" />
                <ENTRY entrytime="00:02:49.25" eventid="1841" heatid="4781" lane="2" />
                <ENTRY entrytime="00:01:16.30" eventid="1992" heatid="4856" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Ludwig" gender="M" lastname="Freutsmiedl" nation="GER" license="263873" athleteid="2603">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.59" eventid="1749" heatid="4680" lane="3" />
                <ENTRY entrytime="00:00:28.65" eventid="1806" heatid="4743" lane="1" />
                <ENTRY entrytime="00:02:15.47" eventid="1820" heatid="4753" lane="5" />
                <ENTRY entrytime="00:02:11.64" eventid="1848" heatid="4791" lane="2" />
                <ENTRY entrytime="00:00:56.44" eventid="1971" heatid="4820" lane="5" />
                <ENTRY entrytime="00:01:01.41" eventid="2013" heatid="4872" lane="5" />
                <ENTRY entrytime="00:04:19.25" eventid="2075" heatid="4910" lane="6" />
                <ENTRY entrytime="00:00:28.63" eventid="2103" heatid="4940" lane="3" />
                <ENTRY entrytime="00:00:27.91" eventid="1912" heatid="5417" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.84" eventid="1961" heatid="4792" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lena" gender="F" lastname="Köhnke" nation="GER" license="284272" athleteid="2612">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.85" eventid="1756" heatid="4689" lane="5" />
                <ENTRY entrytime="00:02:53.20" eventid="1841" heatid="4780" lane="4" />
                <ENTRY entrytime="00:01:19.46" eventid="1992" heatid="4852" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Jana" gender="F" lastname="Lakner" nation="GER" license="281157" athleteid="2616">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.38" eventid="1059" heatid="4666" lane="5" />
                <ENTRY entrytime="00:01:12.97" eventid="1799" heatid="4731" lane="6" />
                <ENTRY entrytime="00:00:31.85" eventid="1855" heatid="4795" lane="6" />
                <ENTRY entrytime="00:00:33.67" eventid="2034" heatid="4885" lane="6" />
                <ENTRY entrytime="00:00:28.45" eventid="2082" heatid="4919" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lukas" gender="M" lastname="Mirsch" nation="GER" license="237415" athleteid="2622">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.80" eventid="1749" heatid="4683" lane="1" />
                <ENTRY entrytime="00:00:57.04" eventid="1778" heatid="4716" lane="4" />
                <ENTRY entrytime="00:00:27.25" eventid="1806" heatid="4743" lane="4" />
                <ENTRY entrytime="00:00:24.65" eventid="1834" heatid="4774" lane="3" />
                <ENTRY entrytime="00:00:53.82" eventid="1971" heatid="4824" lane="3" />
                <ENTRY entrytime="00:02:06.87" eventid="2041" heatid="4894" lane="4" />
                <ENTRY entrytime="00:00:26.28" eventid="2103" heatid="4946" lane="5" />
                <ENTRY entrytime="00:00:27.62" eventid="1912" heatid="4744" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.73" eventid="1898" heatid="4717" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Toni" gender="M" lastname="Schmid" nation="GER" license="227470" athleteid="2630">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.51" eventid="1763" heatid="4703" lane="5" />
                <ENTRY entrytime="00:00:29.57" eventid="1806" heatid="4740" lane="5" />
                <ENTRY entrytime="00:00:25.37" eventid="1834" heatid="4772" lane="5" />
                <ENTRY entrytime="00:00:29.07" eventid="1985" heatid="4848" lane="4" />
                <ENTRY entrytime="00:01:00.70" eventid="2027" heatid="4880" lane="2" />
                <ENTRY entrytime="00:00:27.18" eventid="2103" heatid="4944" lane="4" />
                <ENTRY entrytime="00:01:05.00" eventid="1884" heatid="5368" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Daniel" gender="M" lastname="Siminenko" nation="GER" license="300185" athleteid="2637">
              <ENTRIES>
                <ENTRY entrytime="00:02:11.30" eventid="1749" status="DNS" heatid="4676" lane="2" />
                <ENTRY entrytime="00:01:13.58" eventid="1763" status="DNS" heatid="4697" lane="6" />
                <ENTRY entrytime="00:02:25.22" eventid="1820" status="DNS" heatid="4750" lane="5" />
                <ENTRY entrytime="00:00:27.28" eventid="1834" status="DNS" heatid="4766" lane="3" />
                <ENTRY entrytime="00:00:34.03" eventid="1985" heatid="4841" lane="2" />
                <ENTRY entrytime="00:02:39.38" eventid="2089" heatid="4925" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Tobias" gender="M" lastname="Ulbrich" nation="GER" license="247315" athleteid="2644">
              <ENTRIES>
                <ENTRY entrytime="00:02:08.41" eventid="1749" heatid="4677" lane="3" />
                <ENTRY entrytime="00:02:25.37" eventid="1820" heatid="4750" lane="1" />
                <ENTRY entrytime="00:02:25.12" eventid="1848" heatid="4786" lane="5" />
                <ENTRY entrytime="00:05:08.07" eventid="1999" heatid="4859" lane="2" />
                <ENTRY entrytime="00:04:32.53" eventid="2075" heatid="4908" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4286" nation="GER" region="02" clubid="3328" name="SC DELPHIN Ingolstadt">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Rafaela" gender="F" lastname="Averbeck" nation="GER" license="295302" athleteid="3332">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.60" eventid="1059" heatid="4665" lane="2" />
                <ENTRY entrytime="00:04:40.00" eventid="1827" heatid="4762" lane="4" />
                <ENTRY entrytime="00:19:16.71" eventid="1905" status="RJC">
                  <MEETINFO qualificationtime="00:19:16.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.00" eventid="1978" heatid="4834" lane="3" />
                <ENTRY entrytime="00:09:56.68" eventid="2020" heatid="4875" lane="1">
                  <MEETINFO qualificationtime="00:09:56.68" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Daniel" gender="M" lastname="Chen" nation="GER" license="280055" athleteid="3338">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.60" eventid="1971" heatid="4817" lane="5" />
                <ENTRY entrytime="00:01:06.40" eventid="2013" heatid="4869" lane="1" />
                <ENTRY entrytime="00:00:28.40" eventid="2103" heatid="4941" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Jonas" gender="M" lastname="Drieling" nation="GER" license="280053" athleteid="3345">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.80" eventid="1778" heatid="4713" lane="2" />
                <ENTRY entrytime="00:00:28.40" eventid="1806" heatid="4742" lane="5" />
                <ENTRY entrytime="00:00:25.60" eventid="1834" heatid="4771" lane="2" />
                <ENTRY entrytime="00:00:55.40" eventid="1971" heatid="4822" lane="1" />
                <ENTRY entrytime="00:01:03.40" eventid="2027" heatid="4880" lane="6" />
                <ENTRY entrytime="00:00:26.90" eventid="2103" heatid="4945" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Olivia" gender="F" lastname="Gerrard" nation="GER" license="266868" athleteid="3352">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.10" eventid="1059" heatid="4669" lane="2" />
                <ENTRY entrytime="00:01:07.80" eventid="1785" heatid="4722" lane="1" />
                <ENTRY entrytime="00:00:29.80" eventid="1855" heatid="4800" lane="1" />
                <ENTRY entrytime="00:01:08.80" eventid="2006" heatid="4864" lane="4" />
                <ENTRY entrytime="00:02:31.20" eventid="2055" heatid="4904" lane="6" />
                <ENTRY entrytime="00:02:26.80" eventid="2096" heatid="4937" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Simon" gender="M" lastname="Göpffarth" nation="GER" license="316788" athleteid="3359">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.60" eventid="1749" heatid="4677" lane="5" />
                <ENTRY entrytime="00:00:26.90" eventid="1834" heatid="4767" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Fabian" gender="M" lastname="Heinemann" nation="GER" license="313851" athleteid="3362">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.80" eventid="1778" heatid="4710" lane="6" />
                <ENTRY entrytime="00:00:30.00" eventid="1806" heatid="4740" lane="6" />
                <ENTRY entrytime="00:00:26.00" eventid="1834" heatid="4770" lane="6" />
                <ENTRY entrytime="00:00:56.40" eventid="1971" heatid="4820" lane="2" />
                <ENTRY entrytime="00:01:04.20" eventid="2027" heatid="4878" lane="2" />
                <ENTRY entrytime="00:00:28.00" eventid="2103" heatid="4942" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Larissa" gender="F" lastname="Heinemann" nation="GER" license="313844" athleteid="3369">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.00" eventid="1059" heatid="4667" lane="1" />
                <ENTRY entrytime="00:01:11.80" eventid="1799" heatid="4733" lane="3" />
                <ENTRY entrytime="00:00:31.60" eventid="1855" heatid="4795" lane="3" />
                <ENTRY entrytime="00:01:19.90" eventid="1992" heatid="4852" lane="1" />
                <ENTRY entrytime="00:00:28.40" eventid="2082" heatid="4920" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Joshua" gender="M" lastname="Hollweck" nation="GER" license="313850" athleteid="3375">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.20" eventid="1778" heatid="4712" lane="3" />
                <ENTRY entrytime="00:02:15.60" eventid="1820" heatid="4753" lane="1" />
                <ENTRY entrytime="00:00:55.20" eventid="1971" heatid="4822" lane="2" />
                <ENTRY entrytime="00:02:16.40" eventid="2041" heatid="4893" lane="1" />
                <ENTRY entrytime="00:00:28.10" eventid="2103" heatid="4942" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Iberle" nation="GER" license="313842" athleteid="3381">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.20" eventid="1059" heatid="4664" lane="6" />
                <ENTRY entrytime="00:04:54.00" eventid="1827" heatid="4759" lane="3" />
                <ENTRY entrytime="00:02:20.80" eventid="1978" heatid="4829" lane="4" />
                <ENTRY entrytime="00:02:38.20" eventid="2055" heatid="4898" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lina" gender="F" lastname="Kapfer" nation="GER" license="322567" athleteid="3386">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.60" eventid="1799" heatid="4729" lane="1" />
                <ENTRY entrytime="00:02:54.80" eventid="1841" heatid="4780" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Maria" gender="F" lastname="Kapfer" nation="GER" license="322566" athleteid="3389">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.90" eventid="2034" heatid="4884" lane="4" />
                <ENTRY entrytime="00:02:36.40" eventid="2096" heatid="4932" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sara Maria" gender="F" lastname="Krönert" nation="GER" license="339853" athleteid="3392">
              <ENTRIES>
                <ENTRY entrytime="00:02:33.80" eventid="2096" heatid="4933" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Kuhls" nation="GER" license="265730" athleteid="3394">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.40" eventid="1059" heatid="4668" lane="3" />
                <ENTRY entrytime="00:04:52.00" eventid="1827" heatid="4760" lane="5" />
                <ENTRY entrytime="00:02:17.60" eventid="1978" heatid="4832" lane="5" />
                <ENTRY entrytime="00:00:33.40" eventid="2034" heatid="4885" lane="4" />
                <ENTRY entrytime="00:00:28.60" eventid="2082" heatid="4918" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lukas" gender="M" lastname="Meilinger" nation="GER" license="246338" athleteid="3400">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.60" eventid="1834" heatid="4771" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Raphael" gender="M" lastname="Mooser" nation="GER" license="280056" athleteid="3402">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.40" eventid="1763" heatid="4699" lane="1" />
                <ENTRY entrytime="00:02:23.60" eventid="1820" heatid="4750" lane="4" />
                <ENTRY entrytime="00:00:32.80" eventid="1985" heatid="4842" lane="4" />
                <ENTRY entrytime="00:02:31.20" eventid="2089" heatid="4928" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Sascha" gender="M" lastname="Santa" nation="GER" license="279042" athleteid="3407">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.80" eventid="1749" heatid="4682" lane="5" />
                <ENTRY entrytime="00:02:21.80" eventid="1820" heatid="4751" lane="3" />
                <ENTRY entrytime="00:00:55.60" eventid="1971" heatid="4821" lane="2" />
                <ENTRY entrytime="00:04:13.80" eventid="2075" heatid="4910" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Johanna" gender="F" lastname="Schmid" nation="GER" license="266871" athleteid="3412">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.60" eventid="1756" heatid="4691" lane="5" />
                <ENTRY entrytime="00:01:11.60" eventid="1799" heatid="4735" lane="6" />
                <ENTRY entrytime="00:02:50.00" eventid="1841" heatid="4781" lane="5" />
                <ENTRY entrytime="00:01:18.90" eventid="1992" heatid="4853" lane="6" />
                <ENTRY entrytime="00:02:35.40" eventid="2055" heatid="4900" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Vanessa" gender="F" lastname="Waal" nation="GER" license="301334" athleteid="3418">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.40" eventid="1059" heatid="4666" lane="1" />
                <ENTRY entrytime="00:01:12.90" eventid="1799" heatid="4731" lane="5" />
                <ENTRY entrytime="00:02:20.50" eventid="1978" heatid="4830" lane="5" />
                <ENTRY entrytime="00:00:29.40" eventid="2082" heatid="4915" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4292" nation="GER" region="02" clubid="4087" name="SC Prinz Eugen München">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Alexander Philip" gender="M" lastname="Adami" nation="GER" license="297199" swrid="4829107" athleteid="4103">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.19" eventid="1778" heatid="4710" lane="2" />
                <ENTRY entrytime="00:00:58.07" eventid="1971" heatid="4816" lane="6" />
                <ENTRY entrytime="00:00:28.11" eventid="2103" heatid="4941" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Juliana Andrea" gender="F" lastname="Adami" nation="GER" license="297636" swrid="4829108" athleteid="4107">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.18" eventid="1059" heatid="4666" lane="4" />
                <ENTRY entrytime="00:01:13.22" eventid="1799" heatid="4730" lane="2" />
                <ENTRY entrytime="00:00:30.72" eventid="1855" heatid="4798" lane="3" />
                <ENTRY entrytime="00:02:19.76" eventid="1978" heatid="4831" lane="6" />
                <ENTRY entrytime="00:01:09.83" eventid="2006" heatid="4864" lane="2" />
                <ENTRY entrytime="00:02:36.27" eventid="2055" heatid="4899" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Lyubomir" gender="M" lastname="Agov" nation="GER" license="372659" athleteid="4114">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.50" eventid="1763" heatid="4701" lane="3" />
                <ENTRY entrytime="00:00:26.95" eventid="1985" heatid="4848" lane="3" />
                <ENTRY entrytime="00:01:02.84" eventid="1884" heatid="4704" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Markus" gender="M" lastname="Fischer" nation="GER" license="297634" athleteid="4117">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.49" eventid="1749" heatid="4681" lane="1" />
                <ENTRY entrytime="00:02:13.94" eventid="1848" heatid="4790" lane="5" />
                <ENTRY entrytime="00:00:56.86" eventid="1971" heatid="4819" lane="1" />
                <ENTRY entrytime="00:01:02.22" eventid="2013" heatid="4871" lane="1" />
                <ENTRY entrytime="00:04:22.05" eventid="2075" heatid="4909" lane="2" />
                <ENTRY entrytime="00:09:07.54" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:07.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.01" eventid="1961" heatid="5504" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Jasper" gender="M" lastname="Glindemann" nation="GER" license="309671" athleteid="4124">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.94" eventid="1763" heatid="4698" lane="5" />
                <ENTRY entrytime="00:02:27.77" eventid="1820" heatid="4749" lane="4" />
                <ENTRY entrytime="00:00:31.10" eventid="1985" heatid="4845" lane="5" />
                <ENTRY entrytime="00:01:08.56" eventid="2027" heatid="4877" lane="2" />
                <ENTRY entrytime="00:02:36.40" eventid="2089" heatid="4927" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Kevin" gender="M" lastname="Hültner" nation="GER" license="250305" athleteid="4130">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.87" eventid="1763" heatid="4701" lane="6" />
                <ENTRY entrytime="00:00:30.56" eventid="1985" heatid="4847" lane="6" />
                <ENTRY entrytime="00:02:31.29" eventid="2089" heatid="4927" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Laura" gender="F" lastname="Jaeschke" nation="GER" license="326712" athleteid="4134">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.71" eventid="1059" heatid="4663" lane="6" />
                <ENTRY entrytime="00:04:54.84" eventid="1827" heatid="4759" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Patryk" gender="M" lastname="Laszyca" nation="GER" license="290977" athleteid="4137">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.32" eventid="1778" heatid="4716" lane="1" />
                <ENTRY entrytime="00:00:24.93" eventid="1834" heatid="4774" lane="1" />
                <ENTRY entrytime="00:00:53.86" eventid="1971" heatid="4824" lane="4" />
                <ENTRY entrytime="00:01:03.35" eventid="2027" heatid="4881" lane="6" />
                <ENTRY entrytime="00:00:27.31" eventid="2103" heatid="4944" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Hanna" gender="F" lastname="Pfannes" nation="GER" license="301469" athleteid="4143">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.09" eventid="1756" heatid="4689" lane="6" />
                <ENTRY entrytime="00:02:45.14" eventid="1841" heatid="4783" lane="5" />
                <ENTRY entrytime="00:01:16.20" eventid="1992" heatid="4857" lane="1" />
                <ENTRY entrytime="00:00:33.82" eventid="2034" heatid="4884" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Amelie" gender="F" lastname="Zachenhuber" nation="GER" license="304970" athleteid="4148">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.14" eventid="1059" heatid="4671" lane="2" />
                <ENTRY entrytime="00:00:34.57" eventid="1756" heatid="4692" lane="5" />
                <ENTRY entrytime="00:01:08.67" eventid="1785" heatid="4722" lane="6" />
                <ENTRY entrytime="00:01:10.33" eventid="1799" heatid="4734" lane="5" />
                <ENTRY entrytime="00:00:29.32" eventid="1855" heatid="4961" lane="2" />
                <ENTRY entrytime="00:01:16.36" eventid="1992" heatid="4857" lane="6" />
                <ENTRY entrytime="00:01:07.60" eventid="2006" heatid="4865" lane="1" />
                <ENTRY entrytime="00:00:31.85" eventid="2034" heatid="4889" lane="6" />
                <ENTRY entrytime="00:00:27.53" eventid="2082" heatid="4922" lane="2" />
                <ENTRY entrytime="00:00:29.79" eventid="1940" heatid="5517" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.67" eventid="2048" heatid="4805" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4117" number="1" />
                    <RELAYPOSITION athleteid="4114" number="2" />
                    <RELAYPOSITION athleteid="4103" number="3" />
                    <RELAYPOSITION athleteid="4137" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6524" nation="GER" region="02" clubid="2699" name="SC Regensburg">
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Julia Maria" gender="F" lastname="Grasser" nation="GER" license="179987" athleteid="2700">
              <ENTRIES>
                <ENTRY entrytime="00:02:30.00" eventid="1813" heatid="4746" lane="5" />
                <ENTRY entrytime="00:02:14.15" eventid="1978" heatid="4834" lane="4" />
                <ENTRY entrytime="00:01:07.16" eventid="2006" heatid="4867" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Maximilian" gender="M" lastname="Peter" nation="GER" license="228199" athleteid="2704">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.30" eventid="1806" heatid="4740" lane="4" />
                <ENTRY entrytime="00:02:13.67" eventid="1848" heatid="4791" lane="5" />
                <ENTRY entrytime="00:01:02.14" eventid="2013" heatid="4872" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4296" nation="GER" region="02" clubid="3640" name="SC Wfr. München">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Marvin" gender="M" lastname="Christmann" nation="GER" license="248439" athleteid="3656">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.06" eventid="1763" heatid="4699" lane="5" />
                <ENTRY entrytime="00:00:25.13" eventid="1834" heatid="4773" lane="6" />
                <ENTRY entrytime="00:00:31.36" eventid="1985" heatid="4844" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Dominic" gender="M" lastname="Ehinlanwo" nation="GER" license="302032" athleteid="3660">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.99" eventid="1749" heatid="4684" lane="6" />
                <ENTRY entrytime="00:00:25.02" eventid="1834" heatid="4773" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Bruno" gender="M" lastname="Hediger" nation="GER" license="387694" athleteid="3663">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.24" eventid="1778" heatid="4714" lane="5" />
                <ENTRY entrytime="00:02:11.81" eventid="1820" heatid="4754" lane="1" />
                <ENTRY entrytime="00:00:58.10" eventid="1898" heatid="4717" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julius" gender="M" lastname="Hirschberg" nation="GER" license="333024" athleteid="3666">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.02" eventid="1778" heatid="4711" lane="3" />
                <ENTRY entrytime="00:00:25.73" eventid="1834" heatid="4771" lane="6" />
                <ENTRY entrytime="00:00:27.26" eventid="2103" heatid="4944" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Matthias" gender="M" lastname="Killiches" nation="GER" license="73649" athleteid="3670">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.64" eventid="1763" heatid="4700" lane="3" />
                <ENTRY entrytime="00:00:31.09" eventid="1985" heatid="4845" lane="2" />
                <ENTRY entrytime="00:02:28.00" eventid="2089" heatid="4930" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Jörg" gender="M" lastname="Lukashov" nation="GER" license="252298" athleteid="3674">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.59" eventid="1763" heatid="4702" lane="1" />
                <ENTRY entrytime="00:00:24.05" eventid="1834" heatid="4777" lane="1" />
                <ENTRY entrytime="00:00:53.22" eventid="1971" heatid="4825" lane="5" />
                <ENTRY entrytime="00:00:59.00" eventid="2027" heatid="4879" lane="4" />
                <ENTRY entrytime="00:00:25.82" eventid="2103" heatid="4946" lane="2" />
                <ENTRY entrytime="00:00:23.95" eventid="1947" heatid="4778" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Frida" gender="F" lastname="Mayr" nation="GER" license="356519" athleteid="3680">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.57" eventid="1059" heatid="4668" lane="1" />
                <ENTRY entrytime="00:00:31.62" eventid="1855" heatid="4795" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Viola Jasmine" gender="F" lastname="Provost" nation="GER" license="329228" athleteid="3683">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.22" eventid="1059" heatid="4669" lane="1" />
                <ENTRY entrytime="00:00:28.24" eventid="2082" heatid="4921" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Roman" gender="M" lastname="Roelen" nation="GER" license="283816" athleteid="3686">
              <ENTRIES>
                <ENTRY entrytime="00:02:11.19" eventid="1749" heatid="4676" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="1971" heatid="4813" lane="4" />
                <ENTRY entrytime="00:04:38.00" eventid="2075" heatid="4907" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Alexander" gender="M" lastname="Roschlaub" nation="GER" license="140735" athleteid="3690">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.59" eventid="1749" heatid="4682" lane="4" />
                <ENTRY entrytime="00:00:24.50" eventid="1834" heatid="4775" lane="1" />
                <ENTRY entrytime="00:00:53.31" eventid="1971" heatid="4827" lane="1" />
                <ENTRY entrytime="00:00:24.22" eventid="1947" heatid="5478" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Alexandra" gender="F" lastname="Schäffler" nation="GER" license="231075" athleteid="3694">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.90" eventid="1756" heatid="4691" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Manuel" gender="M" lastname="Straßl" nation="GER" license="132560" athleteid="3696">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.23" eventid="1806" heatid="4743" lane="5" />
                <ENTRY entrytime="00:00:24.70" eventid="1834" heatid="4774" lane="4" />
                <ENTRY entrytime="00:00:54.67" eventid="1971" heatid="4823" lane="1" />
                <ENTRY entrytime="00:01:03.02" eventid="2027" heatid="4880" lane="1" />
                <ENTRY entrytime="00:00:27.00" eventid="2103" heatid="4946" lane="6" />
                <ENTRY entrytime="00:00:24.08" eventid="1947" heatid="5478" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.63" eventid="2048" heatid="4805" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3696" number="1" />
                    <RELAYPOSITION athleteid="3670" number="2" />
                    <RELAYPOSITION athleteid="3663" number="3" />
                    <RELAYPOSITION athleteid="3674" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:42.63" eventid="2232" heatid="4811" lane="4" />
                <ENTRY entrytime="00:02:02.63" eventid="2048" heatid="4805" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3690" number="1" />
                    <RELAYPOSITION athleteid="3656" number="2" />
                    <RELAYPOSITION athleteid="3666" number="3" />
                    <RELAYPOSITION athleteid="3660" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4344" nation="GER" region="02" clubid="3263" name="SCHWIMMVEREIN AUGSBURG 1911 e.V." shortname="SCHWIMMVEREIN AUGSBURG 1911 e.">
          <ATHLETES>
            <ATHLETE birthdate="1989-01-01" firstname="Nadine" gender="F" lastname="Bender" nation="GER" license="197915" athleteid="3264">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.50" eventid="1059" heatid="4673" lane="4" />
                <ENTRY entrytime="00:01:05.20" eventid="1785" heatid="4723" lane="2" />
                <ENTRY entrytime="00:02:08.50" eventid="1978" heatid="4837" lane="2" />
                <ENTRY entrytime="00:00:30.60" eventid="2034" heatid="4888" lane="4" />
                <ENTRY entrytime="00:00:27.30" eventid="2082" heatid="4922" lane="4" />
                <ENTRY entrytime="00:00:59.71" eventid="1863" heatid="5317" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.45" eventid="1891" heatid="5391" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Cara" gender="F" lastname="Gallina" nation="GER" license="299199" athleteid="3270">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.82" eventid="1059" heatid="4664" lane="3" />
                <ENTRY entrytime="00:00:31.50" eventid="1855" heatid="4796" lane="1" />
                <ENTRY entrytime="00:02:16.00" eventid="1978" heatid="4833" lane="6" />
                <ENTRY entrytime="00:00:28.51" eventid="2082" heatid="4919" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Matthias" gender="M" lastname="Kopfmüller" nation="GER" license="137031" athleteid="3275">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.50" eventid="1778" heatid="4715" lane="2" />
                <ENTRY entrytime="00:00:23.40" eventid="1834" heatid="4775" lane="4" />
                <ENTRY entrytime="00:00:51.90" eventid="1971" heatid="4827" lane="2" />
                <ENTRY entrytime="00:00:25.90" eventid="2103" heatid="4945" lane="2" />
                <ENTRY entrytime="00:00:24.26" eventid="5443" heatid="5452" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.26" eventid="1947" heatid="5478" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Andreas" gender="M" lastname="Kornes" nation="GER" license="075398" athleteid="3280">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.40" eventid="1985" heatid="4846" lane="4" />
                <ENTRY entrytime="00:02:23.50" eventid="2089" heatid="4928" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Michelle" gender="F" lastname="Lienhart" nation="GER" license="203026" athleteid="3283">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.74" eventid="1059" heatid="4672" lane="4" />
                <ENTRY entrytime="00:01:06.16" eventid="1799" heatid="4734" lane="3" />
                <ENTRY entrytime="00:00:29.44" eventid="1855" heatid="4800" lane="2" />
                <ENTRY entrytime="00:00:59.49" eventid="1863" heatid="4675" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.35" eventid="1940" heatid="4802" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Oliver" gender="M" lastname="Lienhart" nation="GER" license="248518" athleteid="3287">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.49" eventid="1763" heatid="4699" lane="6" />
                <ENTRY entrytime="00:02:19.55" eventid="1848" heatid="4788" lane="6" />
                <ENTRY entrytime="00:00:57.74" eventid="1971" heatid="4817" lane="6" />
                <ENTRY entrytime="00:01:03.68" eventid="2027" heatid="4878" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Leonie" gender="F" lastname="Mathe" nation="GER" license="215384" athleteid="3292">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.90" eventid="1059" heatid="4674" lane="5" />
                <ENTRY entrytime="00:00:34.00" eventid="1756" heatid="4692" lane="2" />
                <ENTRY entrytime="00:02:47.00" eventid="1841" heatid="4784" lane="6" />
                <ENTRY entrytime="00:01:15.50" eventid="1992" heatid="4855" lane="2" />
                <ENTRY entrytime="00:00:27.50" eventid="2082" heatid="4923" lane="2" />
                <ENTRY entrytime="00:00:33.96" eventid="1877" heatid="4695" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.09" eventid="1954" heatid="5491" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Laura" gender="F" lastname="Popp" nation="GER" license="178550" athleteid="3298">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.60" eventid="1756" heatid="4694" lane="2" />
                <ENTRY entrytime="00:01:07.90" eventid="1799" heatid="4735" lane="2" />
                <ENTRY entrytime="00:02:38.20" eventid="1841" heatid="4782" lane="3" />
                <ENTRY entrytime="00:01:12.90" eventid="1992" heatid="4857" lane="4" />
                <ENTRY entrytime="00:02:27.30" eventid="2055" heatid="4902" lane="2" />
                <ENTRY entrytime="00:00:34.36" eventid="1877" heatid="5355" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.92" eventid="1919" heatid="5404" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:40.61" eventid="1954" heatid="4785" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Lea" gender="F" lastname="Preußner" nation="GER" license="282176" athleteid="3304">
              <ENTRIES>
                <ENTRY entrytime="00:05:26.00" eventid="1771" heatid="4707" lane="2" />
                <ENTRY entrytime="00:01:12.89" eventid="1799" heatid="4731" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Paul" gender="M" lastname="Pucknus" nation="GER" license="264470" athleteid="3307">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.10" eventid="1778" heatid="4711" lane="2" />
                <ENTRY entrytime="00:02:22.25" eventid="1848" heatid="4787" lane="6" />
                <ENTRY entrytime="00:00:58.65" eventid="1971" heatid="4815" lane="1" />
                <ENTRY entrytime="00:02:17.06" eventid="2041" heatid="4894" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Matthias" gender="M" lastname="Schwab" nation="GER" license="132395" athleteid="3312">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.70" eventid="1778" heatid="4715" lane="1" />
                <ENTRY entrytime="00:00:30.20" eventid="1985" heatid="4847" lane="1" />
                <ENTRY entrytime="00:00:25.50" eventid="2103" heatid="4947" lane="4" />
                <ENTRY entrytime="00:00:59.07" eventid="1898" heatid="5465" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Denis" gender="M" lastname="Sczesny" nation="GER" license="350186" athleteid="3316">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.67" eventid="1985" heatid="4841" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Oliver" gender="M" lastname="Sczesny" nation="GER" license="330650" athleteid="3318">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.86" eventid="1763" heatid="4702" lane="5" />
                <ENTRY entrytime="00:00:30.26" eventid="1985" heatid="4846" lane="1" />
                <ENTRY entrytime="00:02:23.53" eventid="2089" heatid="4930" lane="5" />
                <ENTRY entrytime="00:01:04.32" eventid="1884" heatid="5368" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Mark" gender="M" lastname="Toprak" nation="GER" license="346434" athleteid="3322">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.44" eventid="1749" heatid="4680" lane="5" />
                <ENTRY entrytime="00:01:02.89" eventid="1778" heatid="4710" lane="4" />
                <ENTRY entrytime="00:00:56.57" eventid="1971" heatid="4820" lane="1" />
                <ENTRY entrytime="00:02:34.84" eventid="2089" heatid="4927" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.00" eventid="2062" heatid="4807" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3264" number="1" />
                    <RELAYPOSITION athleteid="3298" number="2" />
                    <RELAYPOSITION athleteid="3283" number="3" />
                    <RELAYPOSITION athleteid="3292" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6399" nation="GER" region="02" clubid="3208" name="SG - Elsenfeld/Kleinwallstadt">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Stefanie" gender="F" lastname="Göller" nation="GER" license="245438" athleteid="3217">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.66" eventid="1059" heatid="4668" lane="6" />
                <ENTRY entrytime="00:01:11.70" eventid="1785" heatid="4720" lane="6" />
                <ENTRY entrytime="00:01:12.69" eventid="1799" heatid="4731" lane="3" />
                <ENTRY entrytime="00:00:31.42" eventid="1855" heatid="4796" lane="5" />
                <ENTRY entrytime="00:00:33.48" eventid="2034" heatid="4885" lane="5" />
                <ENTRY entrytime="00:00:28.76" eventid="2082" heatid="4918" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Noelle" gender="F" lastname="Ronalter" nation="GER" license="288664" athleteid="3224">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.03" eventid="1059" heatid="4662" lane="2" />
                <ENTRY entrytime="00:01:13.11" eventid="1785" heatid="4718" lane="3" />
                <ENTRY entrytime="00:01:15.49" eventid="1799" heatid="4728" lane="2" />
                <ENTRY entrytime="00:00:34.21" eventid="2034" heatid="4883" lane="3" />
                <ENTRY entrytime="00:00:29.91" eventid="2082" heatid="4914" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5085" nation="GER" region="02" clubid="4172" name="SG Bamberg">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Benedikt" gender="M" lastname="Dörfler" nation="GER" license="169778" athleteid="4173">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.52" eventid="1749" heatid="4680" lane="1" />
                <ENTRY entrytime="00:00:29.26" eventid="1806" heatid="4740" lane="3" />
                <ENTRY entrytime="00:02:18.13" eventid="1848" heatid="4788" lane="4" />
                <ENTRY entrytime="00:00:56.76" eventid="1971" heatid="4819" lane="5" />
                <ENTRY entrytime="00:01:01.77" eventid="2013" heatid="4871" lane="5" />
                <ENTRY entrytime="00:04:23.39" eventid="2075" heatid="4909" lane="1" />
                <ENTRY entrytime="00:00:28.86" eventid="2103" heatid="4940" lane="2" />
                <ENTRY entrytime="00:02:16.16" eventid="1961" heatid="5504" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Nikolas" gender="M" lastname="Häfner" nation="GER" license="196438" athleteid="4181">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.55" eventid="1806" heatid="4741" lane="3" />
                <ENTRY entrytime="00:00:25.03" eventid="1834" heatid="4773" lane="1" />
                <ENTRY entrytime="00:02:05.45" eventid="1848" heatid="4791" lane="3" />
                <ENTRY entrytime="00:00:51.39" eventid="1971" heatid="4826" lane="4" />
                <ENTRY entrytime="00:00:56.10" eventid="2013" heatid="4873" lane="3" />
                <ENTRY entrytime="00:00:26.80" eventid="2103" heatid="4946" lane="1" />
                <ENTRY entrytime="00:00:27.35" eventid="1912" heatid="4744" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.82" eventid="1961" heatid="4792" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Kevin" gender="M" lastname="Kertész" nation="GER" license="391557" athleteid="4188">
              <ENTRIES>
                <ENTRY entrytime="00:02:08.59" eventid="1749" heatid="4677" lane="4" />
                <ENTRY entrytime="00:02:25.45" eventid="1820" heatid="4750" lane="6" />
                <ENTRY entrytime="00:01:00.17" eventid="1971" heatid="4813" lane="6" />
                <ENTRY entrytime="00:04:39.87" eventid="2075" heatid="4906" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Hanna" gender="F" lastname="Krauß" nation="GER" license="145397" athleteid="4193">
              <ENTRIES>
                <ENTRY entrytime="00:05:09.13" eventid="1771" heatid="4708" lane="5" />
                <ENTRY entrytime="00:04:35.42" eventid="1827" heatid="4763" lane="2" />
                <ENTRY entrytime="00:00:30.97" eventid="1855" heatid="4798" lane="6" />
                <ENTRY entrytime="00:02:10.16" eventid="1978" heatid="4838" lane="1" />
                <ENTRY entrytime="00:09:29.29" eventid="2020" heatid="4876" lane="6">
                  <MEETINFO qualificationtime="00:09:29.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Katrin" gender="F" lastname="Krauß" nation="GER" license="162021" athleteid="4199">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.94" eventid="1059" heatid="4673" lane="5" />
                <ENTRY entrytime="00:04:40.06" eventid="1827" heatid="4762" lane="2" />
                <ENTRY entrytime="00:19:11.45" eventid="1905" status="RJC">
                  <MEETINFO qualificationtime="00:19:11.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.67" eventid="1978" heatid="4836" lane="1" />
                <ENTRY entrytime="00:00:27.84" eventid="2082" heatid="4922" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Dorothea" gender="F" lastname="Rupprecht" nation="GER" license="271055" athleteid="4205">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.36" eventid="2082" heatid="4915" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Julia-Sophia" gender="F" lastname="Scheuermann" nation="GER" license="187882" athleteid="4209">
              <ENTRIES>
                <ENTRY entrytime="00:05:34.66" eventid="1771" heatid="4706" lane="1" />
                <ENTRY entrytime="00:19:25.75" eventid="1905" status="RJC">
                  <MEETINFO qualificationtime="00:19:25.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Bastian" gender="M" lastname="Schorr" nation="GER" license="137664" athleteid="4212">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.76" eventid="1749" heatid="4684" lane="3" />
                <ENTRY entrytime="00:00:56.50" eventid="1778" heatid="4715" lane="3" />
                <ENTRY entrytime="00:00:23.65" eventid="1834" heatid="4776" lane="2" />
                <ENTRY entrytime="00:00:51.17" eventid="1971" heatid="4827" lane="4" />
                <ENTRY entrytime="00:00:58.85" eventid="2027" heatid="4879" lane="3" />
                <ENTRY entrytime="00:00:25.49" eventid="2103" heatid="4945" lane="3" />
                <ENTRY entrytime="00:01:56.80" eventid="1870" heatid="5342" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.14" eventid="5369" heatid="5378" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.14" eventid="1898" heatid="5465" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Corina" gender="F" lastname="Schwandner" nation="GER" license="233736" athleteid="4219">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.68" eventid="1059" heatid="4665" lane="5" />
                <ENTRY entrytime="00:02:19.38" eventid="1978" heatid="4831" lane="2" />
                <ENTRY entrytime="00:00:28.96" eventid="2082" heatid="4917" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Martin" gender="M" lastname="Spörlein" nation="GER" license="169787" athleteid="4223">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.36" eventid="1834" heatid="4776" lane="4" />
                <ENTRY entrytime="00:00:54.66" eventid="1971" heatid="4823" lane="5" />
                <ENTRY entrytime="00:00:23.97" eventid="1947" heatid="5478" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Fabienne" gender="F" lastname="Wenske" nation="GER" license="287819" swrid="5195433" athleteid="4226">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.17" eventid="1059" heatid="4664" lane="1" />
                <ENTRY entrytime="00:05:39.70" eventid="1771" heatid="4705" lane="4" />
                <ENTRY entrytime="00:04:45.59" eventid="1827" heatid="4761" lane="4" />
                <ENTRY entrytime="00:18:55.31" eventid="1905" heatid="4803" lane="1">
                  <MEETINFO qualificationtime="00:18:55.31" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.87" eventid="1978" heatid="4832" lane="2" />
                <ENTRY entrytime="00:02:36.18" eventid="2055" heatid="4899" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Simon" gender="M" lastname="Wicht" nation="GER" license="233738" athleteid="4233">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.51" eventid="1778" heatid="4714" lane="4" />
                <ENTRY entrytime="00:00:27.43" eventid="1806" heatid="4742" lane="4" />
                <ENTRY entrytime="00:02:07.97" eventid="1848" heatid="4789" lane="3" />
                <ENTRY entrytime="00:00:58.80" eventid="2013" status="WDR" heatid="4873" lane="4" />
                <ENTRY entrytime="00:02:09.16" eventid="2041" status="WDR" heatid="4893" lane="4" />
                <ENTRY entrytime="00:00:26.59" eventid="2103" status="WDR" heatid="4947" lane="1" />
                <ENTRY entrytime="00:00:27.68" eventid="1912" heatid="4744" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.98" eventid="1898" heatid="5465" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.92" eventid="1961" heatid="4792" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:46.84" eventid="2048" heatid="4806" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4181" number="1" />
                    <RELAYPOSITION athleteid="4233" number="2" />
                    <RELAYPOSITION athleteid="4212" number="3" />
                    <RELAYPOSITION athleteid="4223" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:36.30" eventid="2232" heatid="4812" lane="5" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5095" nation="GER" region="02" clubid="2755" name="SG Frankenhöhe">
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Johannes" gender="M" lastname="Heinz" nation="GER" license="311886" athleteid="2756">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.00" eventid="1763" heatid="4700" lane="2" />
                <ENTRY entrytime="00:00:30.99" eventid="1985" heatid="4845" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5715" nation="GER" region="02" clubid="3423" name="SG Gundelfingen">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-01" firstname="Charlotte" gender="F" lastname="Joas" nation="GER" license="208201" athleteid="3424">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.19" eventid="1756" heatid="4690" lane="2" />
                <ENTRY entrytime="00:01:19.36" eventid="1992" heatid="4852" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Franziska" gender="F" lastname="Joas" nation="GER" license="155298" athleteid="3427">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.88" eventid="1059" heatid="4667" lane="2" />
                <ENTRY entrytime="00:00:35.26" eventid="1756" heatid="4693" lane="6" />
                <ENTRY entrytime="00:01:12.94" eventid="1799" heatid="4731" lane="1" />
                <ENTRY entrytime="00:00:30.74" eventid="1855" heatid="4798" lane="4" />
                <ENTRY entrytime="00:01:18.02" eventid="1992" heatid="4853" lane="3" />
                <ENTRY entrytime="00:00:28.53" eventid="2082" heatid="4919" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5068" nation="GER" region="02" clubid="2406" name="SG Haßberge">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Jonathan" gender="M" lastname="Bischoff" nation="GER" license="260458" athleteid="2407">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.67" eventid="1763" heatid="4697" lane="4" />
                <ENTRY entrytime="00:00:26.59" eventid="1834" heatid="4767" lane="3" />
                <ENTRY entrytime="00:00:32.35" eventid="1985" heatid="4843" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6768" nation="GER" region="02" clubid="3796" name="SG Mittelfranken">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Varinka" gender="F" lastname="Albert" nation="GER" license="210745" swrid="4193873" athleteid="3801">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.68" eventid="1785" heatid="4723" lane="4" />
                <ENTRY entrytime="00:00:28.41" eventid="1855" heatid="4961" lane="4" />
                <ENTRY entrytime="00:01:04.14" eventid="2006" heatid="4865" lane="4" />
                <ENTRY entrytime="00:00:29.18" eventid="2034" heatid="4889" lane="3" />
                <ENTRY entrytime="00:00:28.13" eventid="2082" heatid="4923" lane="6" />
                <ENTRY entrytime="00:02:18.88" eventid="2096" heatid="4937" lane="4" />
                <ENTRY entrytime="00:01:06.06" eventid="1891" heatid="5391" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.10" eventid="1940" heatid="5517" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Cindy" gender="F" lastname="Blum" nation="GER" license="291192" athleteid="3808">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.57" eventid="1059" heatid="4671" lane="6" />
                <ENTRY entrytime="00:01:12.40" eventid="1785" heatid="4719" lane="5" />
                <ENTRY entrytime="00:04:46.39" eventid="1827" heatid="4761" lane="2" />
                <ENTRY entrytime="NT" eventid="1905" status="RJC" />
                <ENTRY entrytime="00:02:14.65" eventid="1978" heatid="4834" lane="1" />
                <ENTRY entrytime="00:10:02.72" eventid="2020" heatid="4875" lane="6">
                  <MEETINFO qualificationtime="00:10:02.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.04" eventid="2082" heatid="4922" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Bruno" gender="M" lastname="Budde" nation="GER" license="272165" athleteid="3816">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.87" eventid="1749" heatid="4679" lane="6" />
                <ENTRY entrytime="00:17:44.49" eventid="1792" heatid="4726" lane="4">
                  <MEETINFO qualificationtime="00:17:44.49" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.66" eventid="1820" heatid="4752" lane="2" />
                <ENTRY entrytime="00:04:57.75" eventid="1999" heatid="4861" lane="6" />
                <ENTRY entrytime="00:02:19.25" eventid="2041" heatid="4891" lane="3" />
                <ENTRY entrytime="00:00:27.86" eventid="2103" heatid="4942" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Leon" gender="M" lastname="Dresel" nation="GER" license="260105" athleteid="3823">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.09" eventid="1971" heatid="4813" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Justin-Joy" gender="M" lastname="Dutschke" nation="GER" license="293147" athleteid="3825">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.03" eventid="1763" heatid="4699" lane="2" />
                <ENTRY entrytime="00:02:26.46" eventid="1820" heatid="4749" lane="3" />
                <ENTRY entrytime="00:00:57.93" eventid="1971" heatid="4816" lane="2" />
                <ENTRY entrytime="00:00:32.51" eventid="1985" heatid="4843" lane="5" />
                <ENTRY entrytime="00:02:34.03" eventid="2089" heatid="4927" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Dominique" gender="F" lastname="Freisleben" nation="GER" license="242096" athleteid="3835">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.50" eventid="1059" heatid="4671" lane="1" />
                <ENTRY entrytime="00:04:36.00" eventid="1827" heatid="4763" lane="5" />
                <ENTRY entrytime="00:18:26.63" eventid="1905" heatid="4803" lane="3">
                  <MEETINFO qualificationtime="00:18:26.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.00" eventid="1978" heatid="4835" lane="3" />
                <ENTRY entrytime="00:09:30.00" eventid="2020" heatid="4875" lane="3">
                  <MEETINFO qualificationtime="00:09:30.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.00" eventid="2082" heatid="4921" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Mareike" gender="F" lastname="Förster" nation="GER" license="183768" athleteid="3831">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.22" eventid="1756" heatid="4694" lane="4" />
                <ENTRY entrytime="00:01:06.73" eventid="1799" heatid="4735" lane="4" />
                <ENTRY entrytime="00:02:28.55" eventid="1841" heatid="4783" lane="3" />
                <ENTRY entrytime="00:00:34.16" eventid="1877" heatid="5355" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.41" eventid="1919" heatid="4737" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.44" eventid="1954" heatid="4785" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Selina" gender="F" lastname="Herzog" nation="GER" license="274715" athleteid="3842">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.18" eventid="1756" heatid="4688" lane="4" />
                <ENTRY entrytime="00:02:57.83" eventid="1841" heatid="4779" lane="4" />
                <ENTRY entrytime="00:00:32.03" eventid="1855" heatid="4794" lane="2" />
                <ENTRY entrytime="00:01:22.51" eventid="1992" heatid="4850" lane="5" />
                <ENTRY entrytime="00:01:10.47" eventid="2006" heatid="4864" lane="6" />
                <ENTRY entrytime="00:02:39.35" eventid="2055" heatid="4896" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Benno" gender="M" lastname="Hingler" nation="GER" license="242439" athleteid="3849">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.90" eventid="1763" heatid="4698" lane="2" />
                <ENTRY entrytime="00:00:29.84" eventid="1806" heatid="4740" lane="1" />
                <ENTRY entrytime="00:02:22.23" eventid="1820" heatid="4751" lane="2" />
                <ENTRY entrytime="00:00:26.11" eventid="1834" heatid="4769" lane="4" />
                <ENTRY entrytime="00:00:31.72" eventid="1985" heatid="4844" lane="2" />
                <ENTRY entrytime="00:01:03.02" eventid="2027" heatid="4881" lane="1" />
                <ENTRY entrytime="00:02:37.57" eventid="2089" heatid="4926" lane="2" />
                <ENTRY entrytime="00:00:27.36" eventid="2103" heatid="4944" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Hannah" gender="F" lastname="Hofmockel" nation="GER" license="256656" athleteid="3858">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.10" eventid="1756" heatid="4694" lane="5" />
                <ENTRY entrytime="00:01:08.43" eventid="1799" heatid="4734" lane="2" />
                <ENTRY entrytime="00:02:39.01" eventid="1841" heatid="4783" lane="4" />
                <ENTRY entrytime="00:19:09.96" eventid="1905" status="RJC">
                  <MEETINFO qualificationtime="00:19:09.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.65" eventid="1992" heatid="4855" lane="4" />
                <ENTRY entrytime="NT" eventid="2020" status="RJC" />
                <ENTRY entrytime="00:01:09.48" eventid="1919" heatid="4737" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Simon" gender="M" lastname="Jonscher" nation="GER" license="271097" athleteid="3865">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.83" eventid="1749" heatid="4682" lane="1" />
                <ENTRY entrytime="00:01:01.66" eventid="1778" heatid="4712" lane="1" />
                <ENTRY entrytime="00:00:26.00" eventid="1834" heatid="4770" lane="1" />
                <ENTRY entrytime="00:00:55.47" eventid="1971" heatid="4822" lane="6" />
                <ENTRY entrytime="00:01:04.54" eventid="2013" heatid="4870" lane="6" />
                <ENTRY entrytime="00:00:28.23" eventid="2103" heatid="4941" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Jens" gender="M" lastname="Jüttner" nation="GER" license="179877" athleteid="3872">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.59" eventid="1834" heatid="4771" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Daniela" gender="F" lastname="Karst" nation="GER" license="156320" athleteid="3874">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.11" eventid="1756" status="DNS" heatid="4692" lane="3" />
                <ENTRY entrytime="00:01:06.41" eventid="1799" status="DNS" heatid="4736" lane="4" />
                <ENTRY entrytime="00:02:17.97" eventid="1813" status="DNS" heatid="4746" lane="3" />
                <ENTRY entrytime="00:00:28.42" eventid="1855" status="DNS" heatid="4801" lane="4" />
                <ENTRY entrytime="00:01:11.57" eventid="1992" heatid="4857" lane="3" />
                <ENTRY entrytime="00:01:03.15" eventid="2006" heatid="4866" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Kai" gender="M" lastname="Kisberi" nation="GER" license="196491" athleteid="3881">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.15" eventid="1749" heatid="4681" lane="3" />
                <ENTRY entrytime="00:00:26.15" eventid="1834" heatid="4769" lane="2" />
                <ENTRY entrytime="00:00:56.74" eventid="1971" heatid="4819" lane="2" />
                <ENTRY entrytime="00:04:20.97" eventid="2075" heatid="4909" lane="3" />
                <ENTRY entrytime="NT" eventid="2168" status="RJC" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Daniel" gender="M" lastname="Knorr" nation="GER" license="270253" athleteid="3887">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.39" eventid="1778" heatid="4710" lane="5" />
                <ENTRY entrytime="00:02:21.51" eventid="1820" heatid="4752" lane="6" />
                <ENTRY entrytime="00:02:15.36" eventid="1848" heatid="4791" lane="6" />
                <ENTRY entrytime="00:00:57.61" eventid="1971" heatid="4817" lane="1" />
                <ENTRY entrytime="00:01:03.50" eventid="2013" heatid="4870" lane="4" />
                <ENTRY entrytime="00:02:16.82" eventid="2041" heatid="4892" lane="1" />
                <ENTRY entrytime="00:00:28.92" eventid="2103" heatid="4940" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Arthur" gender="M" lastname="Kraft" nation="GER" license="260249" athleteid="3895">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.79" eventid="1971" heatid="4816" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Oliver" gender="M" lastname="Kreißel" nation="GER" license="313677" athleteid="3897">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.71" eventid="1763" heatid="4696" lane="2" />
                <ENTRY entrytime="00:00:33.20" eventid="1985" heatid="4842" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Denis" gender="M" lastname="Kremer" nation="GER" license="302575" athleteid="3900">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.51" eventid="1778" heatid="4709" lane="2" />
                <ENTRY entrytime="00:00:29.10" eventid="1806" heatid="4743" lane="6" />
                <ENTRY entrytime="00:00:26.33" eventid="1834" heatid="4768" lane="3" />
                <ENTRY entrytime="00:02:19.44" eventid="1848" heatid="4788" lane="1" />
                <ENTRY entrytime="00:00:59.48" eventid="1971" heatid="4814" lane="2" />
                <ENTRY entrytime="00:01:04.05" eventid="2013" heatid="4870" lane="5" />
                <ENTRY entrytime="00:01:05.93" eventid="2027" heatid="4877" lane="3" />
                <ENTRY entrytime="00:00:27.03" eventid="2103" heatid="4945" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Elija" gender="M" lastname="Krewer" nation="GER" license="253067" athleteid="3909">
              <ENTRIES>
                <ENTRY entrytime="00:04:36.49" eventid="2075" heatid="4907" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Liv" gender="F" lastname="Krumme" nation="GER" license="281732" athleteid="3911">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.68" eventid="1059" heatid="4670" lane="4" />
                <ENTRY entrytime="00:01:08.91" eventid="1785" heatid="4721" lane="4" />
                <ENTRY entrytime="00:02:15.44" eventid="1978" heatid="4833" lane="2" />
                <ENTRY entrytime="00:00:32.77" eventid="2034" heatid="4886" lane="5" />
                <ENTRY entrytime="00:02:35.02" eventid="2055" heatid="4900" lane="2" />
                <ENTRY entrytime="00:00:28.93" eventid="2082" heatid="4917" lane="3" />
                <ENTRY entrytime="00:02:25.59" eventid="2096" heatid="4935" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Kellie" gender="F" lastname="Messel" nation="GER" license="321746" athleteid="3919">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.75" eventid="1059" heatid="4665" lane="6" />
                <ENTRY entrytime="00:00:38.03" eventid="1756" heatid="4687" lane="6" />
                <ENTRY entrytime="00:04:54.40" eventid="1827" heatid="4759" lane="4" />
                <ENTRY entrytime="00:02:53.89" eventid="1841" heatid="4780" lane="5" />
                <ENTRY entrytime="00:01:20.61" eventid="1992" heatid="4851" lane="1" />
                <ENTRY entrytime="00:02:40.27" eventid="2055" heatid="4896" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Michelle" gender="F" lastname="Messel" nation="GER" license="196996" athleteid="3926">
              <ENTRIES>
                <ENTRY entrytime="00:02:18.23" eventid="1813" heatid="4745" lane="3" />
                <ENTRY entrytime="00:00:28.23" eventid="1855" heatid="4800" lane="3" />
                <ENTRY entrytime="00:01:03.50" eventid="2006" heatid="4865" lane="3" />
                <ENTRY entrytime="00:00:31.80" eventid="2034" heatid="4887" lane="1" />
                <ENTRY entrytime="00:02:22.83" eventid="1933" heatid="4748" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.89" eventid="1940" heatid="4802" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Christoph" gender="M" lastname="Mooser" nation="GER" license="240870" athleteid="3931">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.37" eventid="1763" heatid="4701" lane="1" />
                <ENTRY entrytime="00:00:28.05" eventid="1806" heatid="4741" lane="2" />
                <ENTRY entrytime="00:02:11.16" eventid="1820" heatid="4756" lane="1" />
                <ENTRY entrytime="00:02:14.00" eventid="1848" heatid="4789" lane="5" />
                <ENTRY entrytime="00:00:30.09" eventid="1985" heatid="4848" lane="1" />
                <ENTRY entrytime="00:01:00.21" eventid="2013" heatid="4871" lane="4" />
                <ENTRY entrytime="00:02:23.26" eventid="2089" heatid="4929" lane="2" />
                <ENTRY entrytime="00:00:28.22" eventid="1912" heatid="5417" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.80" eventid="1961" heatid="5504" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Jonas" gender="M" lastname="Mursak" nation="GER" license="196445" athleteid="3939">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.50" eventid="1763" heatid="4703" lane="1" />
                <ENTRY entrytime="00:02:10.00" eventid="1820" heatid="4754" lane="2" />
                <ENTRY entrytime="00:00:30.43" eventid="1985" heatid="4848" lane="6" />
                <ENTRY entrytime="00:00:59.94" eventid="2027" heatid="4881" lane="2" />
                <ENTRY entrytime="00:02:22.50" eventid="2089" heatid="4930" lane="2" />
                <ENTRY entrytime="00:01:05.14" eventid="1884" heatid="5368" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lisa" gender="F" lastname="Mursak" nation="GER" license="196457" athleteid="3945">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.50" eventid="1785" heatid="4723" lane="3" />
                <ENTRY entrytime="00:00:31.03" eventid="1855" heatid="4797" lane="2" />
                <ENTRY entrytime="00:00:29.90" eventid="2034" heatid="4888" lane="3" />
                <ENTRY entrytime="00:02:18.00" eventid="2096" heatid="4935" lane="3" />
                <ENTRY entrytime="00:01:04.72" eventid="1891" heatid="4725" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Katja" gender="F" lastname="Neousypin" nation="GER" license="281139" athleteid="3950">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.63" eventid="1756" heatid="4694" lane="1" />
                <ENTRY entrytime="00:05:34.59" eventid="1771" heatid="4706" lane="5" />
                <ENTRY entrytime="00:02:45.00" eventid="1841" heatid="4784" lane="5" />
                <ENTRY entrytime="00:00:31.41" eventid="1855" heatid="4796" lane="2" />
                <ENTRY entrytime="00:01:15.40" eventid="1992" heatid="4857" lane="2" />
                <ENTRY entrytime="00:01:10.46" eventid="2006" heatid="4864" lane="1" />
                <ENTRY entrytime="00:02:33.79" eventid="2055" heatid="4901" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Tanja" gender="F" lastname="Neubert" nation="GER" license="274074" athleteid="3958">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.43" eventid="1756" heatid="4690" lane="1" />
                <ENTRY entrytime="00:02:45.36" eventid="1841" heatid="4784" lane="1" />
                <ENTRY entrytime="00:01:16.84" eventid="1992" heatid="4856" lane="6" />
                <ENTRY entrytime="00:02:38.75" eventid="2055" heatid="4897" lane="4" />
                <ENTRY entrytime="00:02:46.10" eventid="1954" heatid="5491" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Daniela" gender="F" lastname="Neubig" nation="GER" license="169855" athleteid="3963">
              <ENTRIES>
                <ENTRY entrytime="00:04:59.00" eventid="1771" heatid="4708" lane="4" />
                <ENTRY entrytime="00:02:42.00" eventid="1841" heatid="4784" lane="2" />
                <ENTRY entrytime="00:01:15.77" eventid="1992" heatid="4857" lane="5" />
                <ENTRY entrytime="00:02:23.50" eventid="2055" heatid="4904" lane="2" />
                <ENTRY entrytime="00:02:19.50" eventid="2096" heatid="4936" lane="4" />
                <ENTRY entrytime="00:02:44.11" eventid="1954" heatid="5491" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Jeremias" gender="M" lastname="Pock" nation="GER" license="269306" athleteid="3969">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.77" eventid="1763" heatid="4696" lane="5" />
                <ENTRY entrytime="00:02:22.40" eventid="1820" heatid="4751" lane="6" />
                <ENTRY entrytime="00:02:22.52" eventid="1848" heatid="4786" lane="3" />
                <ENTRY entrytime="00:00:34.35" eventid="1985" heatid="4841" lane="5" />
                <ENTRY entrytime="00:05:05.35" eventid="1999" heatid="4859" lane="3" />
                <ENTRY entrytime="00:02:38.86" eventid="2089" heatid="4926" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Cosima" gender="F" lastname="Rau" nation="GER" license="295229" athleteid="3976">
              <ENTRIES>
                <ENTRY entrytime="00:05:27.81" eventid="1771" heatid="4707" lane="1" />
                <ENTRY entrytime="00:03:06.13" eventid="1841" heatid="4779" lane="1" />
                <ENTRY entrytime="00:01:18.88" eventid="1992" heatid="4853" lane="1" />
                <ENTRY entrytime="00:02:44.43" eventid="2055" heatid="4896" lane="6" />
                <ENTRY entrytime="00:02:41.48" eventid="1954" heatid="5491" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Andreas" gender="M" lastname="Rein" nation="GER" license="278278" athleteid="3981">
              <ENTRIES>
                <ENTRY entrytime="00:01:55.91" eventid="1749" heatid="4683" lane="5" />
                <ENTRY entrytime="00:00:23.47" eventid="1834" heatid="4777" lane="2" />
                <ENTRY entrytime="00:02:09.80" eventid="1848" heatid="4790" lane="4" />
                <ENTRY entrytime="00:00:51.11" eventid="1971" heatid="4826" lane="3" />
                <ENTRY entrytime="00:01:02.43" eventid="2013" heatid="4872" lane="6" />
                <ENTRY entrytime="00:00:25.54" eventid="2103" heatid="4945" lane="4" />
                <ENTRY entrytime="00:00:24.12" eventid="1947" heatid="5478" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Ferdinand" gender="M" lastname="Reng" nation="GER" license="188193" athleteid="3988">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.25" eventid="1834" heatid="4777" lane="4" />
                <ENTRY entrytime="00:00:53.39" eventid="1971" heatid="4826" lane="1" />
                <ENTRY entrytime="00:00:26.22" eventid="2103" heatid="4947" lane="5" />
                <ENTRY entrytime="00:00:23.61" eventid="1947" heatid="4778" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Julian" gender="M" lastname="Richter" nation="GER" license="166195" athleteid="3992">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.87" eventid="1778" heatid="4714" lane="2" />
                <ENTRY entrytime="00:02:10.84" eventid="2041" heatid="4892" lane="2" />
                <ENTRY entrytime="00:00:27.61" eventid="2103" heatid="4943" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Nikita" gender="M" lastname="Rodenko" nation="GER" license="361022" athleteid="3996">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.13" eventid="1749" heatid="4684" lane="1" />
                <ENTRY entrytime="00:02:08.40" eventid="1820" heatid="4756" lane="2" />
                <ENTRY entrytime="00:00:51.15" eventid="1971" heatid="4825" lane="3" />
                <ENTRY entrytime="00:02:12.90" eventid="2041" heatid="4893" lane="5" />
                <ENTRY entrytime="00:08:33.44" eventid="2168" heatid="4809" lane="6">
                  <MEETINFO qualificationtime="00:08:33.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.00" eventid="1870" heatid="4686" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.76" eventid="1926" heatid="5442" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Nele" gender="F" lastname="Rudolph" nation="GER" license="274362" athleteid="4002">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.90" eventid="1059" heatid="4662" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Leonie" gender="F" lastname="Sauer" nation="GER" license="289750" athleteid="4004">
              <ENTRIES>
                <ENTRY entrytime="00:05:29.96" eventid="1771" heatid="4706" lane="4" />
                <ENTRY entrytime="00:02:57.73" eventid="1841" heatid="4779" lane="3" />
                <ENTRY entrytime="00:00:31.94" eventid="1855" heatid="4794" lane="3" />
                <ENTRY entrytime="00:01:21.17" eventid="1992" heatid="4851" lane="6" />
                <ENTRY entrytime="00:02:32.69" eventid="2055" heatid="4901" lane="3" />
                <ENTRY entrytime="00:00:30.08" eventid="2082" heatid="4913" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Helene" gender="F" lastname="Schall" nation="GER" license="309209" athleteid="4011">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.82" eventid="1785" heatid="4721" lane="5" />
                <ENTRY entrytime="00:01:12.29" eventid="1799" heatid="4732" lane="2" />
                <ENTRY entrytime="00:02:20.60" eventid="1978" heatid="4829" lane="3" />
                <ENTRY entrytime="00:00:31.02" eventid="2034" heatid="4889" lane="5" />
                <ENTRY entrytime="00:02:32.04" eventid="2096" heatid="4934" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Ronja" gender="F" lastname="Scharnweber" nation="GER" license="312797" athleteid="4017">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.04" eventid="2082" heatid="4913" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Lars" gender="M" lastname="Schuseil" nation="GER" license="287319" athleteid="4949">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.44" eventid="1749" heatid="4676" lane="3" />
                <ENTRY entrytime="00:00:59.90" eventid="1971" heatid="4813" lane="3" />
                <ENTRY entrytime="00:04:37.87" eventid="2075" heatid="4907" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Alexander" gender="M" lastname="Sinn" nation="GER" license="169871" athleteid="4019">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.73" eventid="1763" heatid="4700" lane="4" />
                <ENTRY entrytime="00:00:25.50" eventid="1834" heatid="4772" lane="6" />
                <ENTRY entrytime="00:00:31.00" eventid="1985" heatid="4845" lane="4" />
                <ENTRY entrytime="00:02:26.87" eventid="2089" heatid="4930" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Anna Lena" gender="F" lastname="Sinn" nation="GER" license="169870" athleteid="4024">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.38" eventid="1756" heatid="4693" lane="4" />
                <ENTRY entrytime="00:00:33.67" eventid="1877" heatid="4695" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Laura" gender="F" lastname="Steuerl" nation="GER" license="316690" athleteid="4953">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.50" eventid="1059" heatid="4668" lane="2" />
                <ENTRY entrytime="00:02:39.13" eventid="1813" heatid="4745" lane="1" />
                <ENTRY entrytime="00:00:32.77" eventid="1855" heatid="4793" lane="2" />
                <ENTRY entrytime="00:19:26.64" eventid="1905" status="RJC">
                  <MEETINFO qualificationtime="00:19:26.64" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.39" eventid="1978" heatid="4833" lane="4" />
                <ENTRY entrytime="NT" eventid="2020" status="RJC" />
                <ENTRY entrytime="00:00:29.28" eventid="2082" heatid="4916" lane="1" />
                <ENTRY entrytime="00:02:35.72" eventid="1933" heatid="5429" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lorenz" gender="M" lastname="Streicher" nation="GER" license="252860" athleteid="4026">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.34" eventid="1749" heatid="4678" lane="5" />
                <ENTRY entrytime="00:01:05.11" eventid="1778" heatid="4709" lane="1" />
                <ENTRY entrytime="00:02:24.62" eventid="1820" heatid="4750" lane="2" />
                <ENTRY entrytime="00:02:21.67" eventid="1848" heatid="4787" lane="5" />
                <ENTRY entrytime="00:05:02.57" eventid="1999" heatid="4860" lane="5" />
                <ENTRY entrytime="00:04:37.27" eventid="2075" heatid="4907" lane="2" />
                <ENTRY entrytime="00:00:29.11" eventid="2103" heatid="4939" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Elena" gender="F" lastname="Tröger" nation="GER" license="307156" athleteid="4034">
              <ENTRIES>
                <ENTRY entrytime="00:02:18.13" eventid="1978" heatid="4832" lane="6" />
                <ENTRY entrytime="00:02:35.10" eventid="2055" heatid="4900" lane="1" />
                <ENTRY entrytime="00:00:29.98" eventid="2082" heatid="4913" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Felicia" gender="F" lastname="Tröger" nation="GER" license="309284" athleteid="4041">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.84" eventid="1756" heatid="4689" lane="4" />
                <ENTRY entrytime="00:01:11.82" eventid="1785" heatid="4719" lane="3" />
                <ENTRY entrytime="00:01:11.56" eventid="1799" heatid="4736" lane="6" />
                <ENTRY entrytime="00:02:53.58" eventid="1841" heatid="4780" lane="2" />
                <ENTRY entrytime="00:00:30.71" eventid="1855" heatid="4799" lane="6" />
                <ENTRY entrytime="00:01:18.79" eventid="1992" heatid="4853" lane="5" />
                <ENTRY entrytime="00:00:34.49" eventid="2034" heatid="4883" lane="2" />
                <ENTRY entrytime="00:02:39.11" eventid="2055" heatid="4897" lane="5" />
                <ENTRY entrytime="00:01:09.93" eventid="1919" heatid="5404" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Emma" gender="F" lastname="Veit" nation="GER" license="301073" athleteid="4050">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.14" eventid="1059" heatid="4667" lane="6" />
                <ENTRY entrytime="00:01:11.10" eventid="1785" heatid="4720" lane="2" />
                <ENTRY entrytime="00:01:10.96" eventid="2006" heatid="4863" lane="4" />
                <ENTRY entrytime="00:02:39.17" eventid="2055" heatid="4897" lane="1" />
                <ENTRY entrytime="00:00:29.46" eventid="2082" heatid="4915" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Karla" gender="F" lastname="Völcker" nation="GER" license="216926" athleteid="4056">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.12" eventid="1059" heatid="4669" lane="5" />
                <ENTRY entrytime="00:01:05.00" eventid="1785" heatid="4724" lane="2" />
                <ENTRY entrytime="00:00:30.93" eventid="1855" heatid="4798" lane="1" />
                <ENTRY entrytime="00:02:15.22" eventid="1978" heatid="4833" lane="3" />
                <ENTRY entrytime="00:00:30.77" eventid="2034" heatid="4887" lane="4" />
                <ENTRY entrytime="00:00:28.48" eventid="2082" heatid="4919" lane="2" />
                <ENTRY entrytime="00:02:21.86" eventid="2096" heatid="4935" lane="2" />
                <ENTRY entrytime="00:01:05.86" eventid="1891" heatid="4725" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Annalena" gender="F" lastname="Wagner" nation="GER" license="297332" athleteid="4064">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.81" eventid="1059" heatid="4672" lane="2" />
                <ENTRY entrytime="00:01:05.98" eventid="1785" heatid="4722" lane="5" />
                <ENTRY entrytime="00:04:39.59" eventid="1827" heatid="4763" lane="6" />
                <ENTRY entrytime="00:02:13.46" eventid="1978" heatid="4835" lane="6" />
                <ENTRY entrytime="00:00:31.44" eventid="2034" heatid="4887" lane="5" />
                <ENTRY entrytime="00:02:19.84" eventid="2096" heatid="4935" lane="4" />
                <ENTRY entrytime="00:00:59.50" eventid="1863" heatid="4675" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.42" eventid="1891" heatid="4725" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Rebecca" gender="F" lastname="Walther" nation="GER" license="292203" athleteid="4071">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.96" eventid="1756" heatid="4687" lane="1" />
                <ENTRY entrytime="00:02:58.72" eventid="1841" heatid="4779" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Deborah" gender="F" lastname="Weber" nation="GER" license="227778" athleteid="4074">
              <ENTRIES>
                <ENTRY entrytime="00:02:25.69" eventid="1813" heatid="4746" lane="2" />
                <ENTRY entrytime="00:00:30.83" eventid="1855" heatid="4798" lane="5" />
                <ENTRY entrytime="NT" eventid="1905" status="RJC" />
                <ENTRY entrytime="00:01:07.13" eventid="2006" heatid="4865" lane="5" />
                <ENTRY entrytime="00:02:25.35" eventid="1933" heatid="4748" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Josefina" gender="F" lastname="Wiesbeck" nation="GER" license="301078" athleteid="4079">
              <ENTRIES>
                <ENTRY entrytime="00:02:29.24" eventid="1813" heatid="4747" lane="5" />
                <ENTRY entrytime="00:00:31.67" eventid="1855" heatid="4795" lane="2" />
                <ENTRY entrytime="00:01:08.16" eventid="2006" heatid="4866" lane="6" />
                <ENTRY entrytime="00:02:25.06" eventid="1933" heatid="4748" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:46.00" eventid="2048" heatid="4806" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3931" number="1" />
                    <RELAYPOSITION athleteid="3939" number="2" />
                    <RELAYPOSITION athleteid="3996" number="3" />
                    <RELAYPOSITION athleteid="3988" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:35.00" eventid="2232" heatid="4812" lane="2" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.00" eventid="2062" heatid="4807" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3945" number="1" />
                    <RELAYPOSITION athleteid="4024" number="2" />
                    <RELAYPOSITION athleteid="3926" number="3" />
                    <RELAYPOSITION athleteid="4064" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:50.00" eventid="2224" heatid="4810" lane="2" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5541" nation="GER" region="02" clubid="2503" name="SG Nordoberpfalz">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Kathrin" gender="F" lastname="Bachmeier" nation="GER" license="262269" athleteid="2504">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.38" eventid="1059" heatid="4669" lane="6" />
                <ENTRY entrytime="00:00:37.81" eventid="1756" heatid="4687" lane="5" />
                <ENTRY entrytime="00:01:13.82" eventid="1785" heatid="4718" lane="5" />
                <ENTRY entrytime="00:01:13.04" eventid="1799" heatid="4730" lane="4" />
                <ENTRY entrytime="00:04:51.69" eventid="1827" heatid="4760" lane="2" />
                <ENTRY entrytime="00:02:19.46" eventid="1978" heatid="4831" lane="1" />
                <ENTRY entrytime="00:02:39.19" eventid="2055" heatid="4897" lane="6" />
                <ENTRY entrytime="00:00:29.16" eventid="2082" heatid="4916" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lukas" gender="M" lastname="Bachmeier" nation="GER" license="210544" athleteid="2513">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.59" eventid="1763" heatid="4698" lane="1" />
                <ENTRY entrytime="00:02:21.85" eventid="1820" heatid="4751" lane="4" />
                <ENTRY entrytime="00:00:32.73" eventid="1985" heatid="4843" lane="6" />
                <ENTRY entrytime="00:02:36.66" eventid="2089" heatid="4926" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Viktoria" gender="F" lastname="Bogner" nation="GER" license="287903" athleteid="2518">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.42" eventid="1059" heatid="4666" lane="6" />
                <ENTRY entrytime="00:00:37.54" eventid="1756" heatid="4687" lane="3" />
                <ENTRY entrytime="00:01:14.66" eventid="1799" heatid="4729" lane="6" />
                <ENTRY entrytime="00:02:20.52" eventid="1978" heatid="4830" lane="1" />
                <ENTRY entrytime="00:01:20.41" eventid="1992" heatid="4851" lane="4" />
                <ENTRY entrytime="00:00:29.74" eventid="2082" heatid="4914" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4305" nation="GER" region="02" clubid="3458" name="SG Oberland T.-I.-P. Penzberg">
          <ATHLETES>
            <ATHLETE birthdate="1990-01-01" firstname="Florian" gender="M" lastname="De Witte" nation="GER" license="307167" athleteid="3459">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.49" eventid="1749" heatid="4679" lane="3" />
                <ENTRY entrytime="00:01:01.20" eventid="1778" heatid="4712" lane="2" />
                <ENTRY entrytime="00:02:15.83" eventid="2041" heatid="4894" lane="1" />
                <ENTRY entrytime="00:00:27.53" eventid="2103" heatid="4943" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Manuel" gender="M" lastname="Genster" nation="GER" license="240652" athleteid="3464">
              <ENTRIES>
                <ENTRY entrytime="00:01:55.88" eventid="1749" heatid="4684" lane="5" />
                <ENTRY entrytime="00:00:55.62" eventid="1778" heatid="4716" lane="3" />
                <ENTRY entrytime="00:00:24.05" eventid="1834" heatid="4775" lane="5" />
                <ENTRY entrytime="00:00:53.15" eventid="1971" heatid="4826" lane="5" />
                <ENTRY entrytime="00:00:25.41" eventid="2103" heatid="4946" lane="3" />
                <ENTRY entrytime="00:00:56.69" eventid="1898" heatid="4717" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Jakob" gender="M" lastname="Hoehler" nation="GER" license="246021" athleteid="3470">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.60" eventid="1763" heatid="4698" lane="3" />
                <ENTRY entrytime="00:00:32.24" eventid="1985" heatid="4843" lane="3" />
                <ENTRY entrytime="00:02:35.80" eventid="2089" heatid="4927" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Philipp" gender="M" lastname="Kirchner" nation="GER" license="131299" athleteid="3474">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.87" eventid="1806" heatid="4743" lane="2" />
                <ENTRY entrytime="00:02:10.00" eventid="1848" heatid="4789" lane="4" />
                <ENTRY entrytime="00:00:58.65" eventid="2013" heatid="4871" lane="3" />
                <ENTRY entrytime="00:00:27.69" eventid="1912" heatid="5417" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Martina Edda" gender="F" lastname="Lickel" nation="GER" license="284991" athleteid="3478">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.97" eventid="1059" heatid="4671" lane="3" />
                <ENTRY entrytime="00:01:08.14" eventid="1785" heatid="4723" lane="6" />
                <ENTRY entrytime="00:02:14.37" eventid="1978" heatid="4834" lane="5" />
                <ENTRY entrytime="00:00:32.21" eventid="2034" heatid="4887" lane="6" />
                <ENTRY entrytime="00:00:27.82" eventid="2082" heatid="4923" lane="5" />
                <ENTRY entrytime="00:01:00.56" eventid="1863" heatid="5317" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Jonathan" gender="M" lastname="Schottenheim" nation="GER" license="306550" athleteid="3484">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.88" eventid="1763" heatid="4697" lane="2" />
                <ENTRY entrytime="00:00:32.33" eventid="1985" heatid="4843" lane="4" />
                <ENTRY entrytime="00:02:38.72" eventid="2089" heatid="4926" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Sebastian" gender="M" lastname="Sonnenstuhl" nation="GER" license="226790" athleteid="3488">
              <ENTRIES>
                <ENTRY entrytime="00:02:17.23" eventid="1820" heatid="4752" lane="3" />
                <ENTRY entrytime="00:00:25.03" eventid="1834" heatid="4773" lane="5" />
                <ENTRY entrytime="00:00:56.22" eventid="1971" heatid="4820" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.00" eventid="2048" heatid="4806" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3474" number="1" />
                    <RELAYPOSITION athleteid="3470" number="2" />
                    <RELAYPOSITION athleteid="3464" number="3" />
                    <RELAYPOSITION athleteid="3488" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6621" nation="GER" region="02" clubid="4242" name="SG Rödental">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Selina" gender="F" lastname="Jenke" nation="GER" license="265832" athleteid="4250">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.85" eventid="1059" heatid="4672" lane="6" />
                <ENTRY entrytime="00:00:30.77" eventid="1855" heatid="4798" lane="2" />
                <ENTRY entrytime="00:00:32.88" eventid="2034" heatid="4886" lane="1" />
                <ENTRY entrytime="00:00:27.70" eventid="2082" heatid="4921" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Danielle" gender="F" lastname="Schuller" nation="GER" license="183972" athleteid="4255">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.43" eventid="1756" heatid="4691" lane="3" />
                <ENTRY entrytime="00:01:11.24" eventid="1799" heatid="4735" lane="1" />
                <ENTRY entrytime="00:01:15.48" eventid="1992" heatid="4856" lane="2" />
                <ENTRY entrytime="00:00:28.59" eventid="2082" heatid="4918" lane="3" />
                <ENTRY entrytime="00:00:34.54" eventid="1877" heatid="5355" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.02" eventid="1919" heatid="5404" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Maike" gender="F" lastname="Schuller" nation="GER" license="183954" athleteid="4260">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.32" eventid="1059" heatid="4663" lane="3" />
                <ENTRY entrytime="00:04:52.31" eventid="1827" heatid="4760" lane="1" />
                <ENTRY entrytime="00:02:20.57" eventid="1978" heatid="4830" lane="6" />
                <ENTRY entrytime="00:02:38.11" eventid="2055" heatid="4898" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.00" eventid="2224" heatid="4810" lane="6" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6423" nation="GER" region="02" clubid="2906" name="SG Stadtwerke München">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Sara" gender="F" lastname="Aringsmann" nation="GER" license="305291" athleteid="2922">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.88" eventid="1059" heatid="4667" lane="4" />
                <ENTRY entrytime="00:00:34.69" eventid="1756" heatid="4693" lane="1" />
                <ENTRY entrytime="00:02:45.21" eventid="1841" heatid="4782" lane="5" />
                <ENTRY entrytime="00:01:16.31" eventid="1992" heatid="4855" lane="1" />
                <ENTRY entrytime="00:02:31.62" eventid="2055" heatid="4903" lane="6" />
                <ENTRY entrytime="00:00:34.09" eventid="1877" heatid="5355" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.32" eventid="1954" heatid="4785" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Yael" gender="M" lastname="Balz" nation="GER" license="318639" athleteid="2928">
              <ENTRIES>
                <ENTRY entrytime="00:17:11.80" eventid="1792" heatid="4726" lane="3" />
                <ENTRY entrytime="00:02:28.30" eventid="1820" heatid="4749" lane="2" />
                <ENTRY entrytime="00:04:15.37" eventid="2075" heatid="4910" lane="5" />
                <ENTRY entrytime="00:08:45.30" eventid="2168" heatid="4808" lane="5">
                  <MEETINFO qualificationtime="00:08:45.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Johanna" gender="F" lastname="Bander" nation="GER" license="281505" athleteid="2933">
              <ENTRIES>
                <ENTRY entrytime="00:04:49.51" eventid="1827" heatid="4760" lane="3" />
                <ENTRY entrytime="00:00:31.74" eventid="1855" heatid="4795" lane="5" />
                <ENTRY entrytime="00:01:22.21" eventid="1992" heatid="4850" lane="3" />
                <ENTRY entrytime="00:02:35.43" eventid="2055" heatid="4899" lane="3" />
                <ENTRY entrytime="00:00:29.07" eventid="2082" heatid="4916" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Janina" gender="F" lastname="Banse" nation="GER" license="234213" athleteid="2939">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.41" eventid="1059" heatid="4674" lane="4" />
                <ENTRY entrytime="00:02:17.80" eventid="1813" heatid="4747" lane="3" />
                <ENTRY entrytime="00:04:22.03" eventid="1827" heatid="4764" lane="4" />
                <ENTRY entrytime="00:02:06.12" eventid="1978" heatid="4838" lane="4" />
                <ENTRY entrytime="00:01:04.11" eventid="2006" heatid="4866" lane="4" />
                <ENTRY entrytime="00:00:27.11" eventid="2082" heatid="4921" lane="3" />
                <ENTRY entrytime="00:00:59.15" eventid="1863" heatid="4675" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.36" eventid="1933" heatid="4748" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Pascal" gender="M" lastname="Borchardt" nation="GER" license="287497" athleteid="2951">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.96" eventid="1749" heatid="4680" lane="4" />
                <ENTRY entrytime="00:01:02.09" eventid="1778" heatid="4711" lane="4" />
                <ENTRY entrytime="00:00:25.42" eventid="1834" heatid="4772" lane="1" />
                <ENTRY entrytime="00:00:55.51" eventid="1971" heatid="4821" lane="4" />
                <ENTRY entrytime="00:00:34.00" eventid="1985" heatid="4841" lane="3" />
                <ENTRY entrytime="00:01:08.46" eventid="2027" heatid="4877" lane="4" />
                <ENTRY entrytime="00:00:27.68" eventid="2103" heatid="4943" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Paulina" gender="F" lastname="Böger" nation="GER" license="202939" athleteid="2946">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.55" eventid="1756" heatid="4692" lane="4" />
                <ENTRY entrytime="00:02:40.10" eventid="1841" heatid="4782" lane="4" />
                <ENTRY entrytime="00:01:13.38" eventid="1992" heatid="4856" lane="4" />
                <ENTRY entrytime="00:02:14.15" eventid="2096" heatid="4937" lane="3" />
                <ENTRY entrytime="00:00:33.54" eventid="1877" heatid="4695" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.66" eventid="1954" heatid="4785" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lisa Marie" gender="F" lastname="Börnigen" nation="GER" license="267312" athleteid="2959">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.77" eventid="1059" heatid="4673" lane="6" />
                <ENTRY entrytime="00:05:14.71" eventid="1771" heatid="4708" lane="6" />
                <ENTRY entrytime="00:02:31.32" eventid="1813" heatid="4745" lane="5" />
                <ENTRY entrytime="00:10:07.84" eventid="2020" status="RJC">
                  <MEETINFO qualificationtime="00:10:07.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.13" eventid="2096" heatid="4934" lane="6" />
                <ENTRY entrytime="00:00:59.99" eventid="1863" heatid="5317" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.16" eventid="1933" heatid="5429" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Benjamin" gender="M" lastname="Campbell-James" nation="GER" license="376054" athleteid="2965">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.63" eventid="1778" heatid="4710" lane="1" />
                <ENTRY entrytime="00:02:14.33" eventid="1820" heatid="4753" lane="4" />
                <ENTRY entrytime="00:02:07.23" eventid="1848" heatid="4790" lane="3" />
                <ENTRY entrytime="00:00:55.12" eventid="1971" heatid="4822" lane="3" />
                <ENTRY entrytime="00:01:00.98" eventid="2013" heatid="4873" lane="5" />
                <ENTRY entrytime="00:04:18.09" eventid="2075" heatid="4910" lane="1" />
                <ENTRY entrytime="00:02:07.71" eventid="1961" heatid="4792" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Elena" gender="F" lastname="Czeschner" nation="GER" license="183021" athleteid="2972">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.50" eventid="1059" heatid="4672" lane="3" />
                <ENTRY entrytime="00:00:27.90" eventid="1855" heatid="4801" lane="3" />
                <ENTRY entrytime="00:01:02.00" eventid="2006" heatid="4867" lane="3" />
                <ENTRY entrytime="00:00:26.31" eventid="2082" heatid="4923" lane="3" />
                <ENTRY entrytime="00:00:29.26" eventid="1940" heatid="4802" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Henning" gender="M" lastname="Dörries" nation="GER" license="220261" athleteid="2977">
              <ENTRIES>
                <ENTRY entrytime="00:01:55.69" eventid="1749" heatid="4685" lane="5" />
                <ENTRY entrytime="00:16:06.02" eventid="1792" heatid="4727" lane="4" />
                <ENTRY entrytime="00:00:25.32" eventid="1834" heatid="4772" lane="2" />
                <ENTRY entrytime="00:04:40.51" eventid="1999" heatid="4862" lane="6" />
                <ENTRY entrytime="00:01:03.55" eventid="2027" heatid="4878" lane="3" />
                <ENTRY entrytime="00:04:06.47" eventid="2075" heatid="4911" lane="3" />
                <ENTRY entrytime="00:08:29.14" eventid="2168" heatid="4809" lane="2">
                  <MEETINFO qualificationtime="00:08:29.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Anastasia" gender="F" lastname="Eftimova" nation="GER" license="323701" athleteid="2985">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.07" eventid="1059" heatid="4662" lane="5" />
                <ENTRY entrytime="00:00:37.02" eventid="1756" heatid="4689" lane="1" />
                <ENTRY entrytime="00:02:57.89" eventid="1841" heatid="4779" lane="2" />
                <ENTRY entrytime="00:01:20.04" eventid="1992" heatid="4852" lane="6" />
                <ENTRY entrytime="00:00:29.74" eventid="2082" heatid="4914" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Veronika" gender="F" lastname="Ehrenbauer" nation="GER" license="106748" athleteid="2991">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.85" eventid="1785" heatid="4724" lane="3" />
                <ENTRY entrytime="00:01:02.93" eventid="1799" heatid="4736" lane="3" />
                <ENTRY entrytime="00:00:27.18" eventid="1855" heatid="4961" lane="3" />
                <ENTRY entrytime="00:01:05.48" eventid="1891" heatid="4725" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.24" eventid="1919" heatid="4737" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.08" eventid="1940" heatid="4802" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Konrad" gender="M" lastname="Fleckenstein" nation="GER" license="247730" athleteid="2995">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.39" eventid="1749" heatid="4681" lane="5" />
                <ENTRY entrytime="00:00:57.50" eventid="1778" heatid="4715" lane="4" />
                <ENTRY entrytime="00:00:24.44" eventid="1834" heatid="4776" lane="1" />
                <ENTRY entrytime="00:00:54.33" eventid="1971" heatid="4823" lane="4" />
                <ENTRY entrytime="00:02:10.00" eventid="2041" heatid="4894" lane="2" />
                <ENTRY entrytime="00:00:25.50" eventid="2103" heatid="4946" lane="4" />
                <ENTRY entrytime="00:00:58.92" eventid="1898" heatid="5465" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Rabea" gender="F" lastname="Gärtner" nation="GER" license="316345" athleteid="3002">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.90" eventid="1059" heatid="4662" lane="3" />
                <ENTRY entrytime="00:00:37.39" eventid="1756" heatid="4688" lane="5" />
                <ENTRY entrytime="00:01:14.20" eventid="1799" heatid="4729" lane="3" />
                <ENTRY entrytime="00:02:51.67" eventid="1841" heatid="4781" lane="6" />
                <ENTRY entrytime="00:01:20.08" eventid="1992" heatid="4851" lane="3" />
                <ENTRY entrytime="00:02:40.18" eventid="2055" heatid="4896" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Benno" gender="M" lastname="Hawe" nation="GER" license="68494" athleteid="3009">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.00" eventid="1763" heatid="4702" lane="4" />
                <ENTRY entrytime="00:00:29.54" eventid="1985" heatid="4847" lane="2" />
                <ENTRY entrytime="00:02:15.00" eventid="2089" heatid="4929" lane="3" />
                <ENTRY entrytime="00:01:04.27" eventid="1884" heatid="5368" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Anna" gender="F" lastname="Herbst" nation="GER" license="250303" athleteid="3013">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.82" eventid="1785" heatid="4723" lane="5" />
                <ENTRY entrytime="00:02:28.47" eventid="1813" heatid="4745" lane="2" />
                <ENTRY entrytime="00:00:29.53" eventid="1855" heatid="4961" lane="5" />
                <ENTRY entrytime="00:01:05.00" eventid="2006" heatid="4867" lane="2" />
                <ENTRY entrytime="00:00:31.72" eventid="2034" heatid="4889" lane="1" />
                <ENTRY entrytime="00:02:28.00" eventid="2055" heatid="4904" lane="1" />
                <ENTRY entrytime="00:02:27.29" eventid="2096" heatid="4936" lane="6" />
                <ENTRY entrytime="00:01:06.21" eventid="1891" heatid="5391" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.09" eventid="1940" heatid="5517" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Anastasia" gender="F" lastname="Ismyrli" nation="GER" license="332675" athleteid="3021">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.71" eventid="1756" heatid="4693" lane="3" />
                <ENTRY entrytime="00:02:38.25" eventid="1841" heatid="4784" lane="4" />
                <ENTRY entrytime="00:00:29.89" eventid="1855" heatid="4961" lane="6" />
                <ENTRY entrytime="00:01:11.63" eventid="1992" heatid="4856" lane="3" />
                <ENTRY entrytime="00:01:05.72" eventid="2006" heatid="4865" lane="2" />
                <ENTRY entrytime="00:00:33.33" eventid="1877" heatid="4695" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.17" eventid="1954" heatid="4785" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Sebastian" gender="M" lastname="Koller" nation="GER" license="184756" athleteid="3027">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.26" eventid="1763" heatid="4703" lane="2" />
                <ENTRY entrytime="00:00:29.42" eventid="1985" heatid="4848" lane="2" />
                <ENTRY entrytime="00:02:16.45" eventid="2089" heatid="4928" lane="3" />
                <ENTRY entrytime="00:01:05.19" eventid="1884" heatid="5368" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Stella" gender="F" lastname="Koltermann" nation="GER" license="245421" athleteid="3031">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.87" eventid="1785" status="DNS" heatid="4720" lane="3" />
                <ENTRY entrytime="00:00:31.17" eventid="1855" status="DNS" heatid="4797" lane="6" />
                <ENTRY entrytime="00:02:14.22" eventid="1978" heatid="4834" lane="2" />
                <ENTRY entrytime="00:00:28.28" eventid="2082" heatid="4920" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Victoria" gender="F" lastname="Kothny" nation="GER" license="274693" athleteid="3201">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.50" eventid="1059" heatid="4672" lane="1" />
                <ENTRY entrytime="00:01:05.50" eventid="1785" heatid="4722" lane="2" />
                <ENTRY entrytime="00:04:41.00" eventid="1827" heatid="4762" lane="1" />
                <ENTRY entrytime="00:02:12.50" eventid="1978" heatid="4835" lane="2" />
                <ENTRY entrytime="00:00:30.41" eventid="2034" heatid="4889" lane="4" />
                <ENTRY entrytime="00:02:21.88" eventid="2096" heatid="4937" lane="5" />
                <ENTRY entrytime="00:01:06.31" eventid="1891" heatid="5391" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Robert" gender="M" lastname="Könneker" nation="GER" license="75201" athleteid="3036">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.49" eventid="1806" heatid="4743" lane="3" />
                <ENTRY entrytime="00:00:22.91" eventid="1834" heatid="4776" lane="3" />
                <ENTRY entrytime="00:00:24.96" eventid="1912" heatid="4744" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.31" eventid="1947" heatid="4778" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Amelie" gender="F" lastname="Liesenfeld" nation="GER" license="301144" athleteid="3039">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.23" eventid="1756" heatid="4690" lane="5" />
                <ENTRY entrytime="00:05:39.47" eventid="1771" heatid="4705" lane="3" />
                <ENTRY entrytime="00:01:14.38" eventid="1799" heatid="4729" lane="4" />
                <ENTRY entrytime="00:02:46.90" eventid="1841" heatid="4782" lane="1" />
                <ENTRY entrytime="00:01:17.21" eventid="1992" heatid="4854" lane="2" />
                <ENTRY entrytime="00:02:38.64" eventid="2055" heatid="4897" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Luisa" gender="F" lastname="Liesenfeld" nation="GER" license="297730" athleteid="3046">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.64" eventid="1059" heatid="4663" lane="1" />
                <ENTRY entrytime="00:04:42.94" eventid="1827" heatid="4762" lane="6" />
                <ENTRY entrytime="00:18:42.01" eventid="1905" heatid="4803" lane="4">
                  <MEETINFO qualificationtime="00:18:42.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.10" eventid="1978" heatid="4832" lane="3" />
                <ENTRY entrytime="00:09:48.60" eventid="2020" heatid="4875" lane="2">
                  <MEETINFO qualificationtime="00:09:48.60" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Anna" gender="F" lastname="Metzler" nation="GER" license="278615" athleteid="3058">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.03" eventid="1059" heatid="4674" lane="1" />
                <ENTRY entrytime="00:01:05.80" eventid="1785" heatid="4724" lane="5" />
                <ENTRY entrytime="00:02:44.59" eventid="1841" heatid="4782" lane="2" />
                <ENTRY entrytime="00:02:06.56" eventid="1978" heatid="4837" lane="4" />
                <ENTRY entrytime="00:01:06.36" eventid="2006" heatid="4866" lane="5" />
                <ENTRY entrytime="00:02:22.81" eventid="2055" heatid="4902" lane="4" />
                <ENTRY entrytime="00:02:23.00" eventid="2096" heatid="4936" lane="5" />
                <ENTRY entrytime="00:00:59.37" eventid="1863" heatid="4675" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.04" eventid="1891" heatid="4725" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Andreas" gender="M" lastname="März" nation="GER" license="301258" athleteid="3052">
              <ENTRIES>
                <ENTRY entrytime="00:17:51.18" eventid="1792" heatid="4726" lane="2" />
                <ENTRY entrytime="00:02:15.00" eventid="1848" heatid="4790" lane="1" />
                <ENTRY entrytime="00:04:50.04" eventid="1999" heatid="4861" lane="1" />
                <ENTRY entrytime="00:01:00.90" eventid="2013" heatid="4871" lane="2" />
                <ENTRY entrytime="00:02:40.53" eventid="2089" heatid="4925" lane="4" />
                <ENTRY entrytime="00:02:11.97" eventid="1961" heatid="4792" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Mara" gender="F" lastname="Münsch" nation="GER" license="280574" athleteid="3066">
              <ENTRIES>
                <ENTRY entrytime="00:05:32.07" eventid="1771" heatid="4706" lane="2" />
                <ENTRY entrytime="00:01:15.49" eventid="1799" heatid="4728" lane="5" />
                <ENTRY entrytime="00:04:50.00" eventid="1827" heatid="4760" lane="4" />
                <ENTRY entrytime="00:02:19.98" eventid="1978" heatid="4830" lane="3" />
                <ENTRY entrytime="00:02:38.79" eventid="2055" heatid="4897" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Max" gender="M" lastname="Nowosad" nation="GER" license="170324" athleteid="3072">
              <ENTRIES>
                <ENTRY entrytime="00:01:48.00" eventid="1749" heatid="4685" lane="3" />
                <ENTRY entrytime="00:02:06.00" eventid="1820" heatid="4756" lane="4" />
                <ENTRY entrytime="00:00:51.76" eventid="1971" heatid="4825" lane="4" />
                <ENTRY entrytime="00:02:05.00" eventid="2041" heatid="4893" lane="3" />
                <ENTRY entrytime="00:03:49.00" eventid="2075" heatid="4912" lane="4" />
                <ENTRY entrytime="NT" eventid="2168" status="RJC" />
                <ENTRY entrytime="00:01:51.42" eventid="1870" heatid="4686" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.94" eventid="1926" heatid="4757" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Christopher" gender="M" lastname="Richter" nation="GER" license="278786" athleteid="3079">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.18" eventid="1749" heatid="4683" lane="2" />
                <ENTRY entrytime="00:01:01.48" eventid="1778" heatid="4712" lane="5" />
                <ENTRY entrytime="00:00:25.16" eventid="1834" heatid="4772" lane="3" />
                <ENTRY entrytime="00:00:53.44" eventid="1971" heatid="4825" lane="1" />
                <ENTRY entrytime="00:04:13.87" eventid="2075" heatid="4910" lane="2" />
                <ENTRY entrytime="00:08:40.79" eventid="2168" heatid="4808" lane="2">
                  <MEETINFO qualificationtime="00:08:39.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.86" eventid="1870" heatid="5342" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Felix" gender="M" lastname="Richtsfeld" nation="GER" license="223387" athleteid="3086">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.00" eventid="1749" heatid="4685" lane="1" />
                <ENTRY entrytime="00:02:12.00" eventid="1820" heatid="4756" lane="6" />
                <ENTRY entrytime="00:00:53.54" eventid="1971" heatid="4827" lane="6" />
                <ENTRY entrytime="00:04:03.00" eventid="2075" heatid="4912" lane="1" />
                <ENTRY entrytime="00:08:35.70" eventid="2168" heatid="4808" lane="4">
                  <MEETINFO qualificationtime="00:08:35.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.33" eventid="1870" heatid="4686" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.90" eventid="1926" heatid="5442" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Derik" gender="M" lastname="Rodrigues" nation="GER" license="245161" athleteid="3092">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.60" eventid="1749" heatid="4679" lane="4" />
                <ENTRY entrytime="00:00:59.11" eventid="1778" heatid="4715" lane="5" />
                <ENTRY entrytime="00:02:19.79" eventid="1820" heatid="4752" lane="5" />
                <ENTRY entrytime="00:00:57.00" eventid="1971" heatid="4818" lane="1" />
                <ENTRY entrytime="00:01:01.93" eventid="2013" heatid="4873" lane="1" />
                <ENTRY entrytime="00:02:10.00" eventid="2041" heatid="4892" lane="4" />
                <ENTRY entrytime="00:00:58.88" eventid="1898" heatid="5465" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Aleksandar" gender="M" lastname="Savic" nation="GER" license="292599" athleteid="3099">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.74" eventid="1749" heatid="4679" lane="1" />
                <ENTRY entrytime="00:01:02.48" eventid="1778" heatid="4711" lane="1" />
                <ENTRY entrytime="00:00:25.98" eventid="1834" heatid="4770" lane="5" />
                <ENTRY entrytime="00:00:56.97" eventid="1971" heatid="4818" lane="2" />
                <ENTRY entrytime="00:01:06.50" eventid="2013" heatid="4869" lane="6" />
                <ENTRY entrytime="00:04:24.68" eventid="2075" heatid="4909" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Dajana" gender="F" lastname="Schlegel" nation="GER" license="158544" athleteid="3106">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.83" eventid="1059" heatid="4670" lane="2" />
                <ENTRY entrytime="00:01:05.00" eventid="1785" heatid="4722" lane="4" />
                <ENTRY entrytime="00:04:29.00" eventid="1827" heatid="4764" lane="1" />
                <ENTRY entrytime="00:02:11.00" eventid="1978" heatid="4837" lane="6" />
                <ENTRY entrytime="00:00:31.40" eventid="2034" heatid="4888" lane="5" />
                <ENTRY entrytime="00:02:28.00" eventid="2055" heatid="4903" lane="1" />
                <ENTRY entrytime="00:02:18.00" eventid="2096" heatid="4936" lane="3" />
                <ENTRY entrytime="00:01:03.72" eventid="1891" heatid="4725" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Lisa Ava" gender="F" lastname="Schlüter" nation="GER" license="310203" athleteid="3114">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.24" eventid="1059" heatid="4666" lane="2" />
                <ENTRY entrytime="00:01:13.25" eventid="1785" heatid="4718" lane="2" />
                <ENTRY entrytime="00:19:00.58" eventid="1905" heatid="4803" lane="6">
                  <MEETINFO qualificationtime="00:19:00.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.09" eventid="1978" heatid="4834" lane="6" />
                <ENTRY entrytime="00:10:03.80" eventid="2020" status="RJC">
                  <MEETINFO qualificationtime="00:09:59.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.37" eventid="2096" heatid="4933" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Marc" gender="M" lastname="Schmid" nation="GER" license="186315" athleteid="3127">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.01" eventid="1763" heatid="4701" lane="4" />
                <ENTRY entrytime="00:02:04.60" eventid="1820" heatid="4755" lane="3" />
                <ENTRY entrytime="00:02:09.05" eventid="1848" heatid="4791" lane="4" />
                <ENTRY entrytime="00:04:23.02" eventid="1999" heatid="4862" lane="3" />
                <ENTRY entrytime="00:02:04.67" eventid="2041" heatid="4894" lane="3" />
                <ENTRY entrytime="00:02:17.62" eventid="2089" heatid="4930" lane="4" />
                <ENTRY entrytime="00:01:03.08" eventid="1884" heatid="4704" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.08" eventid="1926" heatid="4757" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1985-01-01" firstname="Christoph" gender="M" lastname="Thade" nation="GER" license="132608" athleteid="3134">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.00" eventid="1749" heatid="4681" lane="4" />
                <ENTRY entrytime="00:00:25.95" eventid="1806" heatid="4742" lane="3" />
                <ENTRY entrytime="00:00:23.08" eventid="1834" heatid="4775" lane="3" />
                <ENTRY entrytime="00:00:52.00" eventid="1971" heatid="4826" lane="2" />
                <ENTRY entrytime="00:00:57.68" eventid="2013" heatid="4872" lane="3" />
                <ENTRY entrytime="00:00:27.88" eventid="1912" heatid="5417" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Titze" nation="GER" license="272986" athleteid="3140">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.56" eventid="1756" heatid="4694" lane="3" />
                <ENTRY entrytime="00:01:04.18" eventid="1785" heatid="4722" lane="3" />
                <ENTRY entrytime="00:01:04.76" eventid="1799" heatid="4735" lane="3" />
                <ENTRY entrytime="00:00:29.74" eventid="1855" heatid="4801" lane="1" />
                <ENTRY entrytime="00:01:12.72" eventid="1992" heatid="4855" lane="3" />
                <ENTRY entrytime="00:00:30.24" eventid="2034" heatid="4887" lane="3" />
                <ENTRY entrytime="00:02:22.39" eventid="2055" heatid="4903" lane="4" />
                <ENTRY entrytime="00:00:32.56" eventid="1877" heatid="4695" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.38" eventid="1919" heatid="4737" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Sarah" gender="F" lastname="Vidic" nation="GER" license="290443" athleteid="3148">
              <ENTRIES>
                <ENTRY entrytime="00:05:28.09" eventid="1771" heatid="4707" lane="6" />
                <ENTRY entrytime="00:01:07.51" eventid="1785" heatid="4723" lane="1" />
                <ENTRY entrytime="00:00:32.32" eventid="2034" heatid="4886" lane="3" />
                <ENTRY entrytime="00:02:32.79" eventid="2055" heatid="4901" lane="4" />
                <ENTRY entrytime="00:02:24.13" eventid="2096" heatid="4937" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Grant" gender="M" lastname="Wasserman" nation="GER" license="374576" athleteid="3154">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.50" eventid="1749" heatid="4681" lane="6" />
                <ENTRY entrytime="00:01:04.14" eventid="1778" heatid="4709" lane="4" />
                <ENTRY entrytime="00:00:28.88" eventid="1806" heatid="4742" lane="1" />
                <ENTRY entrytime="00:00:24.95" eventid="1834" status="DNS" heatid="4773" lane="4" />
                <ENTRY entrytime="00:00:55.50" eventid="1971" heatid="4821" lane="3" />
                <ENTRY entrytime="00:01:02.28" eventid="2013" heatid="4873" lane="6" />
                <ENTRY entrytime="00:04:27.29" eventid="2075" heatid="4908" lane="3" />
                <ENTRY entrytime="00:00:28.11" eventid="2103" heatid="4941" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Sebastian" gender="M" lastname="Wenk" nation="GER" license="182900" athleteid="3163">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.64" eventid="1749" heatid="4682" lane="2" />
                <ENTRY entrytime="00:01:01.09" eventid="1778" heatid="4713" lane="1" />
                <ENTRY entrytime="00:16:30.00" eventid="1792" heatid="4727" lane="5" />
                <ENTRY entrytime="00:02:15.43" eventid="1820" heatid="4753" lane="2" />
                <ENTRY entrytime="00:02:24.29" eventid="1848" heatid="4786" lane="2" />
                <ENTRY entrytime="00:00:56.95" eventid="1971" heatid="4818" lane="3" />
                <ENTRY entrytime="00:04:48.44" eventid="1999" heatid="4861" lane="5" />
                <ENTRY entrytime="00:01:03.32" eventid="2027" heatid="4879" lane="1" />
                <ENTRY entrytime="00:02:11.49" eventid="2041" heatid="4894" lane="5" />
                <ENTRY entrytime="00:04:10.22" eventid="2075" heatid="4911" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Greta Sophie" gender="F" lastname="Westermann" nation="GER" license="274028" athleteid="3174">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.62" eventid="1059" heatid="4670" lane="3" />
                <ENTRY entrytime="00:01:12.52" eventid="1799" heatid="4732" lane="1" />
                <ENTRY entrytime="00:04:39.57" eventid="1827" heatid="4763" lane="1" />
                <ENTRY entrytime="00:18:48.21" eventid="1905" heatid="4803" lane="2">
                  <MEETINFO qualificationtime="00:18:48.21" />
                </ENTRY>
                <ENTRY entrytime="00:09:53.98" eventid="2020" heatid="4875" lane="5">
                  <MEETINFO qualificationtime="00:09:53.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.54" eventid="2055" heatid="4904" lane="5" />
                <ENTRY entrytime="00:00:28.32" eventid="2082" heatid="4920" lane="5" />
                <ENTRY entrytime="00:01:10.20" eventid="1919" heatid="5404" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lea" gender="F" lastname="Winzer" nation="GER" license="316349" athleteid="3182">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.93" eventid="1785" heatid="4719" lane="1" />
                <ENTRY entrytime="00:01:15.02" eventid="1799" heatid="4728" lane="4" />
                <ENTRY entrytime="00:00:32.00" eventid="1855" heatid="4794" lane="4" />
                <ENTRY entrytime="00:00:33.37" eventid="2034" heatid="4885" lane="3" />
                <ENTRY entrytime="00:02:36.02" eventid="2096" heatid="4933" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Simon" gender="M" lastname="Wittner" nation="GER" license="273514" athleteid="3188">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.23" eventid="1820" heatid="4756" lane="5" />
                <ENTRY entrytime="00:02:11.88" eventid="1848" heatid="4790" lane="2" />
                <ENTRY entrytime="00:04:40.02" eventid="1999" heatid="4862" lane="1" />
                <ENTRY entrytime="00:09:13.63" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:13.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.80" eventid="1926" heatid="5442" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.09" eventid="1961" heatid="4792" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Oliver" gender="M" lastname="Zeidler" nation="GER" license="167736" athleteid="3193">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.00" eventid="1749" heatid="4683" lane="3" />
                <ENTRY entrytime="00:00:23.90" eventid="1834" heatid="4777" lane="5" />
                <ENTRY entrytime="00:00:50.80" eventid="1971" heatid="4827" lane="3" />
                <ENTRY entrytime="00:01:55.02" eventid="1870" heatid="5342" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.42" eventid="1947" heatid="4778" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:38.48" eventid="2048" heatid="4806" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3036" number="1" />
                    <RELAYPOSITION athleteid="3009" number="2" />
                    <RELAYPOSITION athleteid="3072" number="3" />
                    <RELAYPOSITION athleteid="3193" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:29.29" eventid="2232" heatid="4812" lane="4" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.67" eventid="2062" heatid="4807" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2991" number="1" />
                    <RELAYPOSITION athleteid="3140" number="2" />
                    <RELAYPOSITION athleteid="2972" number="3" />
                    <RELAYPOSITION athleteid="2939" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:42.08" eventid="2224" heatid="4810" lane="3" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6695" nation="GER" region="02" clubid="3452" name="SSG Coburg">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Jonas" gender="M" lastname="Colli" nation="GER" license="257089" athleteid="3453">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.21" eventid="1985" heatid="4844" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Kristof" gender="M" lastname="Kalocsai" nation="GER" license="350499" athleteid="3455">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.54" eventid="1834" heatid="4768" lane="6" />
                <ENTRY entrytime="00:00:59.66" eventid="1971" heatid="4814" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4330" nation="GER" region="02" clubid="2532" name="SSG Neptun Germering e.V.">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Claudia" gender="F" lastname="Dobmeier" nation="GER" license="299888" athleteid="2586">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.85" eventid="2082" heatid="4914" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Mareike" gender="F" lastname="Feller" nation="GER" license="218202" athleteid="2540">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.23" eventid="1785" heatid="4721" lane="2" />
                <ENTRY entrytime="00:01:12.20" eventid="1799" heatid="4733" lane="6" />
                <ENTRY entrytime="00:00:30.64" eventid="1855" heatid="4799" lane="5" />
                <ENTRY entrytime="00:00:32.20" eventid="2034" heatid="4888" lane="6" />
                <ENTRY entrytime="00:00:28.84" eventid="2082" heatid="4918" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Emily" gender="F" lastname="Gallow" nation="GER" license="384453" athleteid="2593">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.55" eventid="1059" heatid="4663" lane="2" />
                <ENTRY entrytime="00:01:14.57" eventid="1799" heatid="4729" lane="5" />
                <ENTRY entrytime="00:00:31.32" eventid="1855" heatid="4796" lane="4" />
                <ENTRY entrytime="00:00:28.57" eventid="2082" heatid="4919" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Franziska" gender="F" lastname="Godau" nation="GER" license="219095" athleteid="2533">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.37" eventid="2082" heatid="4920" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Miriam" gender="F" lastname="Karcher" nation="GER" license="316822" athleteid="2588">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.62" eventid="1756" heatid="4689" lane="3" />
                <ENTRY entrytime="00:01:22.35" eventid="1992" heatid="4850" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Elisa" gender="F" lastname="Lex" nation="GER" license="323971" athleteid="2591">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.51" eventid="1756" heatid="4688" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Laura" gender="F" lastname="Obermayer" nation="GER" license="280497" athleteid="2560">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.57" eventid="1756" heatid="4691" lane="2" />
                <ENTRY entrytime="00:05:16.03" eventid="1771" heatid="4707" lane="4" />
                <ENTRY entrytime="00:04:43.20" eventid="1827" heatid="4761" lane="3" />
                <ENTRY entrytime="00:02:47.49" eventid="1841" heatid="4783" lane="6" />
                <ENTRY entrytime="00:01:17.49" eventid="1992" heatid="4854" lane="1" />
                <ENTRY entrytime="00:02:27.90" eventid="2055" heatid="4903" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Matthias" gender="M" lastname="Rips" nation="GER" license="226730" athleteid="2546">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.98" eventid="1763" heatid="4697" lane="3" />
                <ENTRY entrytime="00:01:00.28" eventid="1778" heatid="4714" lane="6" />
                <ENTRY entrytime="00:02:18.39" eventid="1820" heatid="4752" lane="4" />
                <ENTRY entrytime="00:00:30.94" eventid="1985" heatid="4846" lane="6" />
                <ENTRY entrytime="00:01:02.64" eventid="2027" heatid="4880" lane="5" />
                <ENTRY entrytime="00:02:29.00" eventid="2089" heatid="4929" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Maximilian" gender="M" lastname="Stadler" nation="GER" license="242037" athleteid="2535">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.49" eventid="1806" heatid="4739" lane="1" />
                <ENTRY entrytime="00:00:27.32" eventid="1834" heatid="4766" lane="2" />
                <ENTRY entrytime="00:02:22.75" eventid="1848" heatid="4786" lane="4" />
                <ENTRY entrytime="00:01:05.68" eventid="2013" heatid="4869" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Nele" gender="F" lastname="Ströbel" nation="GER" license="299265" athleteid="2575">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.95" eventid="1059" heatid="4664" lane="2" />
                <ENTRY entrytime="00:04:54.83" eventid="1827" heatid="4759" lane="2" />
                <ENTRY entrytime="00:00:31.59" eventid="1855" heatid="4796" lane="6" />
                <ENTRY entrytime="00:01:11.06" eventid="2006" heatid="4863" lane="2" />
                <ENTRY entrytime="00:02:37.51" eventid="2055" heatid="4898" lane="3" />
                <ENTRY entrytime="00:00:29.32" eventid="2082" heatid="4916" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Nikita" gender="M" lastname="Tsvetkov" nation="GER" license="265703" athleteid="2582">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.37" eventid="1806" heatid="4738" lane="2" />
                <ENTRY entrytime="00:00:27.29" eventid="1834" heatid="4766" lane="4" />
                <ENTRY entrytime="00:00:59.22" eventid="1971" heatid="4814" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Leopold" gender="M" lastname="Wahl" nation="GER" license="246999" athleteid="2553">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.93" eventid="1778" heatid="4709" lane="3" />
                <ENTRY entrytime="00:00:29.13" eventid="1806" heatid="4742" lane="6" />
                <ENTRY entrytime="00:02:12.74" eventid="1848" heatid="4789" lane="2" />
                <ENTRY entrytime="00:00:56.94" eventid="1971" heatid="4819" lane="6" />
                <ENTRY entrytime="00:01:02.48" eventid="2013" heatid="4871" lane="6" />
                <ENTRY entrytime="00:00:27.97" eventid="2103" heatid="4942" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Maximilian" gender="M" lastname="Wipplinger" nation="GER" license="293163" athleteid="2567">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.11" eventid="1749" heatid="4682" lane="3" />
                <ENTRY entrytime="00:16:36.80" eventid="1792" heatid="4727" lane="1" />
                <ENTRY entrytime="00:02:12.71" eventid="1820" heatid="4755" lane="6" />
                <ENTRY entrytime="00:00:54.23" eventid="1971" heatid="4823" lane="3" />
                <ENTRY entrytime="00:04:38.84" eventid="1999" heatid="4862" lane="5" />
                <ENTRY entrytime="00:01:02.71" eventid="2027" heatid="4879" lane="5" />
                <ENTRY entrytime="00:04:09.87" eventid="2075" heatid="4911" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4331" nation="GER" region="02" clubid="3705" name="SSKC Poseidon Aschaffenburg">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Justin" gender="M" lastname="Arapaj" nation="GER" license="243492" swrid="4613309" athleteid="3712">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.03" eventid="1749" heatid="4678" lane="4" />
                <ENTRY entrytime="00:02:20.45" eventid="1848" heatid="4787" lane="3" />
                <ENTRY entrytime="00:00:55.73" eventid="1971" heatid="4821" lane="1" />
                <ENTRY entrytime="00:01:04.50" eventid="2013" heatid="4870" lane="1" />
                <ENTRY entrytime="00:00:27.98" eventid="2103" heatid="4942" lane="5" />
                <ENTRY entrytime="00:02:16.10" eventid="1961" heatid="5504" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Cäcilia" gender="F" lastname="Bausback" nation="GER" license="308503" athleteid="3718">
              <ENTRIES>
                <ENTRY entrytime="00:05:29.90" eventid="1771" heatid="4706" lane="3" />
                <ENTRY entrytime="00:04:55.89" eventid="1827" heatid="4758" lane="4" />
                <ENTRY entrytime="00:00:32.11" eventid="1855" heatid="4793" lane="3" />
                <ENTRY entrytime="00:18:51.87" eventid="1905" heatid="4803" lane="5">
                  <MEETINFO qualificationtime="00:18:51.87" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.38" eventid="2006" heatid="4864" lane="5" />
                <ENTRY entrytime="00:02:37.59" eventid="2055" heatid="4898" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Lisa" gender="F" lastname="Diener" nation="GER" license="192721" athleteid="3725">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.15" eventid="1059" heatid="4671" lane="5" />
                <ENTRY entrytime="00:00:29.62" eventid="1855" heatid="4800" lane="5" />
                <ENTRY entrytime="00:00:28.26" eventid="2082" heatid="4920" lane="3" />
                <ENTRY entrytime="00:00:30.23" eventid="1940" heatid="5517" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Sebastian" gender="M" lastname="Feser" nation="GER" license="173941" athleteid="3729">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.09" eventid="1778" heatid="4716" lane="6" />
                <ENTRY entrytime="00:00:29.34" eventid="1806" heatid="4740" lane="2" />
                <ENTRY entrytime="00:00:25.28" eventid="1834" heatid="4772" lane="4" />
                <ENTRY entrytime="00:00:55.33" eventid="1971" heatid="4822" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Fabienne" gender="F" lastname="Krüger" nation="GER" license="297473" athleteid="3734">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.00" eventid="1059" heatid="4664" lane="5" />
                <ENTRY entrytime="00:04:48.63" eventid="1827" heatid="4761" lane="1" />
                <ENTRY entrytime="00:19:10.47" eventid="1905" status="RJC">
                  <MEETINFO qualificationtime="00:19:10.47" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.75" eventid="1978" heatid="4833" lane="1" />
                <ENTRY entrytime="00:10:14.45" eventid="2020" status="RJC">
                  <MEETINFO qualificationtime="00:10:14.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.42" eventid="2096" heatid="4932" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Dovlat" gender="M" lastname="Mirzoev" nation="GER" license="297743" athleteid="3741">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.56" eventid="1763" heatid="4697" lane="1" />
                <ENTRY entrytime="00:00:27.40" eventid="1834" heatid="4765" lane="2" />
                <ENTRY entrytime="00:00:58.36" eventid="1971" heatid="4815" lane="2" />
                <ENTRY entrytime="00:00:34.01" eventid="1985" heatid="4841" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Ilyas" gender="M" lastname="Mirzoev" nation="GER" license="297744" athleteid="3746">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.66" eventid="1763" heatid="4696" lane="1" />
                <ENTRY entrytime="00:00:26.81" eventid="1834" heatid="4767" lane="2" />
                <ENTRY entrytime="00:00:57.80" eventid="1971" heatid="4816" lane="4" />
                <ENTRY entrytime="00:00:28.92" eventid="2103" heatid="4939" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Anna" gender="F" lastname="Reibenspiess" nation="GER" license="297472" athleteid="3751">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.40" eventid="1059" heatid="4673" lane="1" />
                <ENTRY entrytime="00:01:10.40" eventid="1785" heatid="4721" lane="6" />
                <ENTRY entrytime="00:04:39.82" eventid="1827" heatid="4762" lane="3" />
                <ENTRY entrytime="00:18:21.28" eventid="1905" heatid="4804" lane="6">
                  <MEETINFO qualificationtime="00:18:21.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.48" eventid="1978" heatid="4837" lane="1" />
                <ENTRY entrytime="00:09:35.39" eventid="2020" heatid="4875" lane="4">
                  <MEETINFO qualificationtime="00:09:35.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.86" eventid="2096" heatid="4934" lane="3" />
                <ENTRY entrytime="00:00:59.81" eventid="1863" heatid="5317" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Niklas" gender="M" lastname="Reibenspiess" nation="GER" license="168669" athleteid="3759">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.70" eventid="1763" heatid="4702" lane="6" />
                <ENTRY entrytime="00:02:11.48" eventid="1820" heatid="4755" lane="1" />
                <ENTRY entrytime="00:02:21.03" eventid="1848" heatid="4787" lane="2" />
                <ENTRY entrytime="00:00:54.08" eventid="1971" heatid="4824" lane="5" />
                <ENTRY entrytime="00:04:47.13" eventid="1999" heatid="4861" lane="2" />
                <ENTRY entrytime="00:02:25.50" eventid="2089" heatid="4928" lane="5" />
                <ENTRY entrytime="00:02:09.83" eventid="1926" heatid="5442" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Hanna" gender="F" lastname="Seubert" nation="GER" license="257093" athleteid="3766">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.43" eventid="1756" heatid="4692" lane="6" />
                <ENTRY entrytime="00:01:11.48" eventid="1785" heatid="4720" lane="5" />
                <ENTRY entrytime="00:02:51.75" eventid="1841" heatid="4780" lane="3" />
                <ENTRY entrytime="00:01:18.39" eventid="1992" heatid="4853" lane="4" />
                <ENTRY entrytime="00:00:33.42" eventid="2034" heatid="4885" lane="2" />
                <ENTRY entrytime="00:00:28.10" eventid="2082" heatid="4921" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Philipp" gender="M" lastname="Walter" nation="GER" license="284784" athleteid="3773">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.85" eventid="1749" heatid="4678" lane="6" />
                <ENTRY entrytime="00:17:51.36" eventid="1792" heatid="4726" lane="5" />
                <ENTRY entrytime="00:00:30.72" eventid="1806" heatid="4739" lane="6" />
                <ENTRY entrytime="00:02:18.98" eventid="1848" heatid="4788" lane="5" />
                <ENTRY entrytime="00:04:58.00" eventid="1999" heatid="4860" lane="3" />
                <ENTRY entrytime="00:04:31.31" eventid="2075" heatid="4908" lane="4" />
                <ENTRY entrytime="00:09:16.88" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:16.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.30" eventid="2048" heatid="4805" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3729" number="1" />
                    <RELAYPOSITION athleteid="3759" number="2" />
                    <RELAYPOSITION athleteid="3746" number="3" />
                    <RELAYPOSITION athleteid="3712" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:42.43" eventid="2232" heatid="4811" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3729" number="1" />
                    <RELAYPOSITION athleteid="3759" number="2" />
                    <RELAYPOSITION athleteid="3712" number="3" />
                    <RELAYPOSITION athleteid="3746" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.20" eventid="2062" heatid="4807" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3751" number="1" />
                    <RELAYPOSITION athleteid="3766" number="2" />
                    <RELAYPOSITION athleteid="3718" number="3" />
                    <RELAYPOSITION athleteid="3725" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:55.78" eventid="2224" heatid="4810" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3725" number="1" />
                    <RELAYPOSITION athleteid="3751" number="2" />
                    <RELAYPOSITION athleteid="3766" number="3" />
                    <RELAYPOSITION athleteid="3734" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4347" nation="GER" region="02" clubid="4572" name="SV Bayreuth">
          <ATHLETES>
            <ATHLETE birthdate="1991-01-01" firstname="Christoph" gender="M" lastname="Argauer" nation="GER" license="134500" athleteid="4573">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.17" eventid="1749" heatid="4680" lane="2" />
                <ENTRY entrytime="00:01:09.96" eventid="1763" heatid="4699" lane="3" />
                <ENTRY entrytime="00:00:56.32" eventid="1971" heatid="4820" lane="4" />
                <ENTRY entrytime="00:00:32.10" eventid="1985" heatid="4844" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Jette" gender="F" lastname="Barthmann" nation="GER" license="297427" athleteid="4578">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.02" eventid="1785" heatid="4719" lane="6" />
                <ENTRY entrytime="00:00:31.21" eventid="1855" heatid="4796" lane="3" />
                <ENTRY entrytime="00:01:10.73" eventid="2006" heatid="4863" lane="3" />
                <ENTRY entrytime="00:00:34.09" eventid="2034" heatid="4884" lane="6" />
                <ENTRY entrytime="00:02:37.31" eventid="2055" heatid="4899" lane="6" />
                <ENTRY entrytime="00:02:36.81" eventid="2096" heatid="4932" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Marc Oliver" gender="M" lastname="Birkle" nation="GER" license="269134" athleteid="4585">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.98" eventid="1749" heatid="4678" lane="3" />
                <ENTRY entrytime="00:00:26.05" eventid="1834" heatid="4769" lane="3" />
                <ENTRY entrytime="00:00:56.95" eventid="1971" heatid="4818" lane="4" />
                <ENTRY entrytime="00:00:32.78" eventid="1985" heatid="4842" lane="3" />
                <ENTRY entrytime="00:04:33.07" eventid="2075" heatid="4908" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1991-01-01" firstname="Maximilian" gender="M" lastname="Deichsel" nation="GER" license="138788" athleteid="4591">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.20" eventid="1778" heatid="4715" lane="6" />
                <ENTRY entrytime="00:02:11.11" eventid="1820" heatid="4754" lane="5" />
                <ENTRY entrytime="00:04:45.15" eventid="1999" heatid="4861" lane="4" />
                <ENTRY entrytime="00:00:59.14" eventid="5369" heatid="5378" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.71" eventid="1926" heatid="5442" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Carmen" gender="F" lastname="Gräbner" nation="GER" license="297780" athleteid="4595">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.85" eventid="1756" heatid="4689" lane="2" />
                <ENTRY entrytime="00:05:27.19" eventid="1771" heatid="4707" lane="5" />
                <ENTRY entrytime="00:02:50.30" eventid="1841" heatid="4781" lane="1" />
                <ENTRY entrytime="00:01:19.50" eventid="1992" heatid="4852" lane="5" />
                <ENTRY entrytime="00:02:33.85" eventid="2055" heatid="4901" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Nico" gender="M" lastname="Heilmann" nation="GER" license="291040" athleteid="4601">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.72" eventid="1985" heatid="4840" lane="3" />
                <ENTRY entrytime="00:02:42.39" eventid="2089" heatid="4925" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Luisa" gender="F" lastname="Kauper" nation="GER" license="305148" athleteid="4604">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.71" eventid="1756" heatid="4687" lane="2" />
                <ENTRY entrytime="00:02:48.42" eventid="1841" heatid="4781" lane="3" />
                <ENTRY entrytime="00:01:20.46" eventid="1992" heatid="4851" lane="2" />
                <ENTRY entrytime="00:02:35.98" eventid="2055" heatid="4899" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Florian" gender="M" lastname="Müller" nation="GER" license="266235" athleteid="4609">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.58" eventid="1763" heatid="4703" lane="6" />
                <ENTRY entrytime="00:01:00.46" eventid="1778" heatid="4713" lane="3" />
                <ENTRY entrytime="00:02:14.13" eventid="1820" heatid="4753" lane="3" />
                <ENTRY entrytime="00:00:55.14" eventid="1971" heatid="4822" lane="4" />
                <ENTRY entrytime="00:00:31.16" eventid="1985" heatid="4845" lane="1" />
                <ENTRY entrytime="00:02:23.81" eventid="2089" heatid="4929" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Selina" gender="F" lastname="Müller" nation="GER" license="242742" athleteid="4616">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.00" eventid="1785" heatid="4724" lane="6" />
                <ENTRY entrytime="00:00:31.77" eventid="2034" heatid="4888" lane="1" />
                <ENTRY entrytime="00:02:24.16" eventid="2096" heatid="4936" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Stefanie" gender="F" lastname="Raps" nation="GER" license="234205" athleteid="4620">
              <ENTRIES>
                <ENTRY entrytime="00:02:34.70" eventid="1813" heatid="4746" lane="1" />
                <ENTRY entrytime="00:04:52.54" eventid="1827" heatid="4760" lane="6" />
                <ENTRY entrytime="00:02:21.48" eventid="1978" heatid="4829" lane="5" />
                <ENTRY entrytime="00:01:11.67" eventid="2006" heatid="4863" lane="5" />
                <ENTRY entrytime="00:02:34.79" eventid="2055" heatid="4900" lane="4" />
                <ENTRY entrytime="00:02:30.37" eventid="1933" heatid="5429" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.00" eventid="2048" heatid="4805" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4591" number="1" />
                    <RELAYPOSITION athleteid="4573" number="2" />
                    <RELAYPOSITION athleteid="4609" number="3" />
                    <RELAYPOSITION athleteid="4585" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:44.00" eventid="2232" heatid="4811" lane="2" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4356" nation="GER" region="02" clubid="2436" name="SV GR.-W. Holzkirchen">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-01" firstname="Ludwig" gender="M" lastname="Huber" nation="GER" license="181978" athleteid="2437">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.00" eventid="1749" heatid="4682" lane="6" />
                <ENTRY entrytime="00:01:10.63" eventid="1763" heatid="4698" lane="4" />
                <ENTRY entrytime="00:01:01.15" eventid="1778" heatid="4713" lane="6" />
                <ENTRY entrytime="00:00:24.54" eventid="1834" heatid="4776" lane="6" />
                <ENTRY entrytime="00:00:54.20" eventid="1971" heatid="4824" lane="6" />
                <ENTRY entrytime="00:00:32.00" eventid="1985" heatid="4844" lane="5" />
                <ENTRY entrytime="00:00:27.26" eventid="2103" heatid="4944" lane="2" />
                <ENTRY entrytime="00:00:24.26" eventid="5443" heatid="5452" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5713" nation="GER" region="02" clubid="2488" name="SV Hengersberg">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Fabian" gender="M" lastname="Miller" nation="GER" license="282389" athleteid="2489">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.08" eventid="1971" heatid="4815" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Erik" gender="M" lastname="Stögbauer" nation="GER" license="291450" athleteid="2491">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.16" eventid="1806" heatid="4738" lane="4" />
                <ENTRY entrytime="00:00:27.00" eventid="1834" heatid="4767" lane="6" />
                <ENTRY entrytime="00:01:00.13" eventid="1971" heatid="4813" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4341" nation="GER" region="02" clubid="4628" name="SV Hof 1911 e. V.">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Leon" gender="M" lastname="Richter" nation="GER" license="270159" athleteid="4636">
              <ENTRIES>
                <ENTRY entrytime="00:18:47.39" eventid="1792" heatid="4726" lane="1" />
                <ENTRY entrytime="00:00:26.95" eventid="1834" heatid="4767" lane="1" />
                <ENTRY entrytime="00:00:59.88" eventid="1971" heatid="4814" lane="6" />
                <ENTRY entrytime="00:04:39.47" eventid="2075" heatid="4906" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Matthias" gender="M" lastname="Schmidt" nation="GER" license="209569" athleteid="4641">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.33" eventid="1834" heatid="4768" lane="4" />
                <ENTRY entrytime="00:00:27.80" eventid="2103" heatid="4942" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4364" nation="GER" region="02" clubid="3247" name="SV Ottobrunn 1970 e.V.">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Birte" gender="F" lastname="Schiemann" nation="GER" license="260141" athleteid="3248">
              <ENTRIES>
                <ENTRY entrytime="00:02:19.40" eventid="1978" heatid="4831" lane="5" />
                <ENTRY entrytime="00:00:33.00" eventid="2034" heatid="4886" lane="6" />
                <ENTRY entrytime="00:00:28.76" eventid="2082" heatid="4918" lane="2" />
                <ENTRY entrytime="00:02:32.49" eventid="2096" heatid="4934" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4384" nation="GER" region="02" clubid="2445" name="SV Wacker Burghausen">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Verena" gender="F" lastname="Bergmann" nation="GER" license="295270" athleteid="2446">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.00" eventid="1785" heatid="4719" lane="4" />
                <ENTRY entrytime="00:01:13.00" eventid="1799" heatid="4730" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Yannick" gender="M" lastname="Buschhardt" nation="GER" license="227101" athleteid="2449">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.00" eventid="1806" heatid="4742" lane="2" />
                <ENTRY entrytime="00:00:24.50" eventid="1834" heatid="4777" lane="6" />
                <ENTRY entrytime="00:00:53.60" eventid="1971" heatid="4825" lane="6" />
                <ENTRY entrytime="00:00:59.00" eventid="2013" heatid="4872" lane="4" />
                <ENTRY entrytime="00:00:27.31" eventid="1912" heatid="4744" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Marina" gender="F" lastname="Hammerl" nation="GER" license="284445" athleteid="2454">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.56" eventid="1059" heatid="4668" lane="5" />
                <ENTRY entrytime="00:02:32.00" eventid="1813" heatid="4747" lane="1" />
                <ENTRY entrytime="00:00:31.00" eventid="1855" heatid="4797" lane="3" />
                <ENTRY entrytime="00:02:16.50" eventid="1978" heatid="4832" lane="4" />
                <ENTRY entrytime="00:01:08.00" eventid="2006" heatid="4867" lane="6" />
                <ENTRY entrytime="00:00:29.50" eventid="2082" heatid="4915" lane="1" />
                <ENTRY entrytime="00:02:29.62" eventid="1933" heatid="5429" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Dominik" gender="M" lastname="Kohlschmid" nation="GER" license="242746" athleteid="2461">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.50" eventid="1763" heatid="4701" lane="5" />
                <ENTRY entrytime="00:00:58.00" eventid="1778" heatid="4716" lane="2" />
                <ENTRY entrytime="00:02:07.00" eventid="1820" heatid="4754" lane="4" />
                <ENTRY entrytime="00:00:54.40" eventid="1971" heatid="4823" lane="2" />
                <ENTRY entrytime="00:00:30.00" eventid="1985" heatid="4846" lane="5" />
                <ENTRY entrytime="00:00:59.00" eventid="2027" heatid="4880" lane="4" />
                <ENTRY entrytime="00:02:27.00" eventid="2089" heatid="4928" lane="1" />
                <ENTRY entrytime="00:00:27.00" eventid="2103" heatid="4947" lane="6" />
                <ENTRY entrytime="00:02:08.00" eventid="1926" heatid="4757" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.05" eventid="1898" heatid="4717" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Paulina" gender="F" lastname="Sandner" nation="GER" license="316586" athleteid="2470">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.50" eventid="1059" heatid="4668" lane="4" />
                <ENTRY entrytime="00:00:35.70" eventid="1756" heatid="4691" lane="1" />
                <ENTRY entrytime="00:01:10.00" eventid="1799" heatid="4735" lane="5" />
                <ENTRY entrytime="00:01:17.00" eventid="1992" heatid="4854" lane="3" />
                <ENTRY entrytime="00:00:29.00" eventid="2082" heatid="4917" lane="1" />
                <ENTRY entrytime="00:01:10.08" eventid="1919" heatid="5404" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Marlene" gender="F" lastname="Sommoggy von" nation="GER" license="304160" athleteid="2476">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.00" eventid="1756" heatid="4690" lane="3" />
                <ENTRY entrytime="00:01:12.00" eventid="1799" heatid="4733" lane="2" />
                <ENTRY entrytime="00:02:48.00" eventid="1841" heatid="4782" lane="6" />
                <ENTRY entrytime="00:01:17.00" eventid="1992" heatid="4854" lane="4" />
                <ENTRY entrytime="00:00:34.18" eventid="1877" heatid="5355" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:44.28" eventid="1954" heatid="5491" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4387" nation="GER" region="02" clubid="4648" name="SV Weiden">
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Lisa" gender="F" lastname="Biersack" nation="GER" license="225273" athleteid="4649">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.57" eventid="1785" heatid="4724" lane="4" />
                <ENTRY entrytime="00:01:10.75" eventid="1799" heatid="4736" lane="1" />
                <ENTRY entrytime="00:00:29.92" eventid="1855" heatid="4800" lane="6" />
                <ENTRY entrytime="00:00:31.02" eventid="2034" heatid="4887" lane="2" />
                <ENTRY entrytime="00:02:23.95" eventid="2096" heatid="4935" lane="5" />
                <ENTRY entrytime="00:01:07.04" eventid="1891" heatid="5391" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Alina" gender="F" lastname="Zimmermann" nation="GER" license="193325" athleteid="4655">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.03" eventid="1059" heatid="4671" lane="4" />
                <ENTRY entrytime="00:01:11.69" eventid="1799" heatid="4734" lane="6" />
                <ENTRY entrytime="00:00:30.49" eventid="1855" heatid="4799" lane="3" />
                <ENTRY entrytime="00:02:12.72" eventid="1978" heatid="4835" lane="5" />
                <ENTRY entrytime="00:01:07.53" eventid="2006" heatid="4866" lane="1" />
                <ENTRY entrytime="00:00:28.03" eventid="2082" heatid="4923" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4339" nation="GER" region="02" clubid="3493" name="SV Würzburg 05">
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Leonie Antonia" gender="F" lastname="Beck" nation="GER" license="186145" athleteid="3502">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.64" eventid="1059" heatid="4674" lane="3" />
                <ENTRY entrytime="00:02:27.87" eventid="1841" heatid="4784" lane="3" />
                <ENTRY entrytime="00:01:57.90" eventid="1978" heatid="4838" lane="3" />
                <ENTRY entrytime="00:02:11.87" eventid="2055" heatid="4904" lane="3" />
                <ENTRY entrytime="00:00:57.46" eventid="1863" heatid="4675" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.07" eventid="1954" heatid="4785" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Maximilian" gender="M" lastname="Beck" nation="GER" license="161820" athleteid="3507">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.46" eventid="1763" heatid="4702" lane="3" />
                <ENTRY entrytime="00:02:03.48" eventid="1820" heatid="4756" lane="3" />
                <ENTRY entrytime="00:00:23.65" eventid="1834" heatid="4775" lane="2" />
                <ENTRY entrytime="00:00:29.13" eventid="1985" heatid="4847" lane="4" />
                <ENTRY entrytime="00:00:57.94" eventid="2027" heatid="4880" lane="3" />
                <ENTRY entrytime="00:01:04.19" eventid="1884" heatid="4704" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.51" eventid="1926" heatid="4757" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Sebastian Aurelius" gender="M" lastname="Beck" nation="GER" license="236295" athleteid="3513">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.28" eventid="1749" heatid="4683" lane="4" />
                <ENTRY entrytime="00:02:06.50" eventid="1820" heatid="4755" lane="4" />
                <ENTRY entrytime="00:00:52.39" eventid="1971" heatid="4825" lane="2" />
                <ENTRY entrytime="00:03:58.67" eventid="2075" heatid="4912" lane="2" />
                <ENTRY entrytime="00:08:30.03" eventid="2168" heatid="4809" lane="1">
                  <MEETINFO qualificationtime="00:08:30.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.95" eventid="1870" heatid="5342" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.63" eventid="1926" heatid="4757" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Max" gender="M" lastname="Brandenstein" nation="GER" license="312913" athleteid="3519">
              <ENTRIES>
                <ENTRY entrytime="00:16:41.28" eventid="1792" heatid="4727" lane="6" />
                <ENTRY entrytime="00:00:26.30" eventid="1834" heatid="4769" lane="6" />
                <ENTRY entrytime="00:00:56.74" eventid="1971" heatid="4819" lane="4" />
                <ENTRY entrytime="00:04:11.51" eventid="2075" heatid="4910" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Frederik" gender="M" lastname="Bär" nation="GER" license="249941" athleteid="3497">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.50" eventid="1806" heatid="4741" lane="5" />
                <ENTRY entrytime="00:00:24.78" eventid="1834" heatid="4774" lane="2" />
                <ENTRY entrytime="00:00:55.00" eventid="1971" heatid="4823" lane="6" />
                <ENTRY entrytime="00:01:02.00" eventid="2027" heatid="4881" lane="5" />
                <ENTRY entrytime="00:00:27.77" eventid="1912" heatid="5417" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Klemens" gender="M" lastname="Degenhardt" nation="GER" license="140643" athleteid="3524">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.79" eventid="1763" heatid="4703" lane="3" />
                <ENTRY entrytime="00:02:14.23" eventid="1848" heatid="4791" lane="1" />
                <ENTRY entrytime="00:00:28.04" eventid="1985" heatid="4847" lane="3" />
                <ENTRY entrytime="00:02:12.26" eventid="2089" heatid="4930" lane="3" />
                <ENTRY entrytime="00:08:34.84" eventid="2168" heatid="4808" lane="3">
                  <MEETINFO qualificationtime="00:08:34.84" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.99" eventid="1884" heatid="4704" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Carolin" gender="F" lastname="Dorfner" nation="GER" license="244045" athleteid="3530">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.60" eventid="1059" heatid="4673" lane="2" />
                <ENTRY entrytime="00:02:19.55" eventid="1813" heatid="4746" lane="4" />
                <ENTRY entrytime="00:00:29.55" eventid="1855" heatid="4801" lane="5" />
                <ENTRY entrytime="00:01:03.53" eventid="2006" heatid="4867" lane="4" />
                <ENTRY entrytime="00:02:21.52" eventid="2055" heatid="4904" lane="4" />
                <ENTRY entrytime="00:00:59.51" eventid="1863" heatid="5317" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.28" eventid="1933" heatid="4748" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Romy" gender="F" lastname="Dreher" nation="GER" license="269748" athleteid="3546">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1059" heatid="4672" lane="5" />
                <ENTRY entrytime="00:04:22.48" eventid="1827" heatid="4764" lane="2" />
                <ENTRY entrytime="00:17:40.54" eventid="1905" heatid="4804" lane="2">
                  <MEETINFO qualificationtime="00:17:40.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.11" eventid="1978" heatid="4836" lane="4" />
                <ENTRY entrytime="00:09:09.01" eventid="2020" heatid="4876" lane="4">
                  <MEETINFO qualificationtime="00:09:09.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.24" eventid="1863" heatid="5317" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Tim" gender="M" lastname="Dreher" nation="GER" license="205376" athleteid="3552">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.16" eventid="1749" heatid="4684" lane="4" />
                <ENTRY entrytime="00:02:10.31" eventid="1820" heatid="4755" lane="5" />
                <ENTRY entrytime="00:02:06.68" eventid="2041" heatid="4892" lane="3" />
                <ENTRY entrytime="00:08:53.45" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:08:53.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.92" eventid="1870" heatid="5342" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Luise" gender="F" lastname="Dörries" nation="GER" license="162166" athleteid="3536">
              <ENTRIES>
                <ENTRY entrytime="00:05:15.89" eventid="1771" heatid="4707" lane="3" />
                <ENTRY entrytime="00:04:31.25" eventid="1827" heatid="4763" lane="3" />
                <ENTRY entrytime="00:17:32.78" eventid="1905" heatid="4804" lane="4">
                  <MEETINFO qualificationtime="00:17:32.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.94" eventid="1978" heatid="4838" lane="6" />
                <ENTRY entrytime="00:09:14.39" eventid="2020" heatid="4876" lane="2">
                  <MEETINFO qualificationtime="00:09:14.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Susanne" gender="F" lastname="Dörries" nation="GER" license="157347" athleteid="3542">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.00" eventid="1978" heatid="4836" lane="6" />
                <ENTRY entrytime="NT" eventid="2020" status="RJC" />
                <ENTRY entrytime="00:02:28.00" eventid="2096" heatid="4935" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Dix" gender="M" lastname="Eisenbraun" nation="GER" license="176717" athleteid="3557">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="1763" heatid="4699" lane="4" />
                <ENTRY entrytime="00:02:14.00" eventid="1820" heatid="4754" lane="6" />
                <ENTRY entrytime="00:02:13.00" eventid="2041" heatid="4892" lane="5" />
                <ENTRY entrytime="00:02:27.00" eventid="2089" heatid="4929" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Sebastian" gender="M" lastname="Greß" nation="GER" license="138833" athleteid="3562">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.00" eventid="1778" heatid="4714" lane="3" />
                <ENTRY entrytime="00:00:24.00" eventid="1834" heatid="4776" lane="5" />
                <ENTRY entrytime="00:00:30.00" eventid="1985" heatid="4847" lane="5" />
                <ENTRY entrytime="00:00:59.00" eventid="2027" heatid="4881" lane="4" />
                <ENTRY entrytime="00:00:25.00" eventid="2103" heatid="4947" lane="3" />
                <ENTRY entrytime="00:00:55.47" eventid="1898" heatid="4717" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.68" eventid="1947" heatid="4778" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lars" gender="M" lastname="Grundheber" nation="GER" license="234237" athleteid="3568">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.89" eventid="1749" heatid="4684" lane="2" />
                <ENTRY entrytime="00:02:05.13" eventid="1820" heatid="4754" lane="3" />
                <ENTRY entrytime="00:04:25.52" eventid="1999" heatid="4862" lane="4" />
                <ENTRY entrytime="00:03:59.65" eventid="2075" heatid="4912" lane="5" />
                <ENTRY entrytime="00:08:29.14" eventid="2168" heatid="4809" lane="5">
                  <MEETINFO qualificationtime="00:08:29.14" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.41" eventid="1870" heatid="4686" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.67" eventid="1926" heatid="4757" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Alina" gender="F" lastname="Hennl" nation="GER" license="173169" athleteid="3574">
              <ENTRIES>
                <ENTRY entrytime="00:04:54.33" eventid="1771" status="DNS" heatid="4708" lane="3" />
                <ENTRY entrytime="00:02:18.46" eventid="1813" status="DNS" heatid="4747" lane="4" />
                <ENTRY entrytime="00:02:09.35" eventid="1978" heatid="4836" lane="2" />
                <ENTRY entrytime="00:02:18.44" eventid="2055" heatid="4902" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Svenja" gender="F" lastname="Herbert" nation="GER" license="304086" athleteid="3579">
              <ENTRIES>
                <ENTRY entrytime="00:05:10.90" eventid="1771" heatid="4708" lane="1" />
                <ENTRY entrytime="00:04:30.00" eventid="1827" heatid="4764" lane="6" />
                <ENTRY entrytime="00:17:55.70" eventid="1905" heatid="4804" lane="1">
                  <MEETINFO qualificationtime="00:17:55.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.00" eventid="1978" heatid="4838" lane="5" />
                <ENTRY entrytime="00:02:27.99" eventid="2055" heatid="4902" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Alina" gender="F" lastname="Jungklaus" nation="GER" license="249937" athleteid="3585">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.81" eventid="1059" heatid="4673" lane="3" />
                <ENTRY entrytime="00:04:07.45" eventid="1827" heatid="4764" lane="3" />
                <ENTRY entrytime="00:16:55.04" eventid="1905" heatid="4804" lane="3">
                  <MEETINFO qualificationtime="00:16:55.04" />
                </ENTRY>
                <ENTRY entrytime="00:01:59.16" eventid="1978" heatid="4837" lane="3" />
                <ENTRY entrytime="00:00:27.11" eventid="2082" heatid="4923" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Lena" gender="F" lastname="Kalla" nation="GER" license="143081" athleteid="3591">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.00" eventid="1799" heatid="4734" lane="4" />
                <ENTRY entrytime="00:00:29.00" eventid="1855" heatid="4800" lane="4" />
                <ENTRY entrytime="00:00:31.00" eventid="2034" heatid="4888" lane="2" />
                <ENTRY entrytime="00:02:20.00" eventid="2096" heatid="4937" lane="2" />
                <ENTRY entrytime="00:01:06.17" eventid="1919" heatid="4737" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.16" eventid="1940" heatid="4802" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Jakob" gender="M" lastname="Markowski" nation="GER" license="154737" athleteid="3596">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.76" eventid="1763" heatid="4703" lane="4" />
                <ENTRY entrytime="00:00:22.86" eventid="1834" heatid="4777" lane="3" />
                <ENTRY entrytime="00:00:28.79" eventid="1985" heatid="4846" lane="3" />
                <ENTRY entrytime="00:00:57.45" eventid="2027" heatid="4881" lane="3" />
                <ENTRY entrytime="00:01:02.39" eventid="1884" heatid="4704" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.47" eventid="1947" heatid="4778" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1990-01-01" firstname="Sören" gender="M" lastname="Meißner" nation="GER" license="106221" athleteid="3601">
              <ENTRIES>
                <ENTRY entrytime="00:07:58.29" eventid="2168" heatid="4809" lane="4">
                  <MEETINFO qualificationtime="00:07:58.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Laura" gender="F" lastname="Neumann" nation="GER" license="249654" athleteid="3603">
              <ENTRIES>
                <ENTRY entrytime="00:05:00.00" eventid="1771" heatid="4708" lane="2" />
                <ENTRY entrytime="00:02:44.00" eventid="1841" heatid="4783" lane="2" />
                <ENTRY entrytime="00:02:10.00" eventid="1978" heatid="4837" lane="5" />
                <ENTRY entrytime="00:02:26.00" eventid="2055" heatid="4903" lane="2" />
                <ENTRY entrytime="00:02:43.04" eventid="1954" heatid="5491" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Leonie" gender="F" lastname="Neumann" nation="GER" license="249655" athleteid="3608">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.56" eventid="1059" heatid="4674" lane="6" />
                <ENTRY entrytime="00:04:32.16" eventid="1827" heatid="4763" lane="4" />
                <ENTRY entrytime="00:17:55.14" eventid="1905" heatid="4804" lane="5">
                  <MEETINFO qualificationtime="00:17:55.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.00" eventid="1978" heatid="4836" lane="5" />
                <ENTRY entrytime="00:09:23.26" eventid="2020" heatid="4876" lane="1">
                  <MEETINFO qualificationtime="00:09:19.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Natalie" gender="F" lastname="Schnabel" nation="GER" license="299453" athleteid="3614">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.69" eventid="1059" heatid="4665" lane="1" />
                <ENTRY entrytime="00:00:37.43" eventid="1756" heatid="4688" lane="1" />
                <ENTRY entrytime="00:02:55.37" eventid="1841" heatid="4780" lane="6" />
                <ENTRY entrytime="00:01:18.78" eventid="1992" heatid="4853" lane="2" />
                <ENTRY entrytime="00:02:35.06" eventid="2055" heatid="4900" lane="5" />
                <ENTRY entrytime="00:00:29.00" eventid="2082" heatid="4917" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Ruwen" gender="M" lastname="Straub" nation="GER" license="148906" athleteid="3621">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.19" eventid="1749" heatid="4685" lane="4" />
                <ENTRY entrytime="00:02:17.32" eventid="1848" heatid="4789" lane="6" />
                <ENTRY entrytime="00:00:52.90" eventid="1971" heatid="4827" lane="5" />
                <ENTRY entrytime="00:03:45.56" eventid="2075" heatid="4912" lane="3" />
                <ENTRY entrytime="00:07:54.96" eventid="2168" heatid="4809" lane="3">
                  <MEETINFO qualificationtime="00:07:54.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.64" eventid="1870" heatid="4686" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Shay" gender="M" lastname="Toledano" nation="GER" license="365525" athleteid="3627">
              <ENTRIES>
                <ENTRY entrytime="00:15:48.48" eventid="1792" heatid="4727" lane="3" />
                <ENTRY entrytime="00:04:45.03" eventid="1999" heatid="4861" lane="3" />
                <ENTRY entrytime="00:04:08.47" eventid="2075" heatid="4911" lane="2" />
                <ENTRY entrytime="00:08:47.66" eventid="2168" heatid="4808" lane="1">
                  <MEETINFO qualificationtime="00:08:47.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Svenja" gender="F" lastname="Zihsler" nation="GER" license="151222" athleteid="3632">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.52" eventid="1978" heatid="4836" lane="3" />
                <ENTRY entrytime="00:08:40.16" eventid="2020" heatid="4876" lane="3">
                  <MEETINFO qualificationtime="00:08:40.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.74" eventid="2055" heatid="4903" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:44.00" eventid="2048" heatid="4806" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3497" number="1" />
                    <RELAYPOSITION athleteid="3524" number="2" />
                    <RELAYPOSITION athleteid="3562" number="3" />
                    <RELAYPOSITION athleteid="3596" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:26.89" eventid="2232" heatid="4812" lane="3" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:01:58.00" eventid="2062" heatid="4807" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3591" number="1" />
                    <RELAYPOSITION athleteid="3502" number="2" />
                    <RELAYPOSITION athleteid="3530" number="3" />
                    <RELAYPOSITION athleteid="3585" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:47.00" eventid="2224" heatid="4810" lane="4" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5806" nation="GER" region="02" clubid="2708" name="Team Buron Kaufbeuren">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Nadja" gender="F" lastname="Amrhein" nation="GER" license="262168" swrid="4491234" athleteid="2709">
              <ENTRIES>
                <ENTRY entrytime="00:01:17.55" eventid="1992" heatid="4854" lane="6" />
                <ENTRY entrytime="00:02:32.52" eventid="2055" heatid="4902" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Katharina" gender="F" lastname="Breunig" nation="GER" license="299621" athleteid="2712">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.64" eventid="1059" heatid="4663" lane="5" />
                <ENTRY entrytime="00:00:37.66" eventid="1756" heatid="4687" lane="4" />
                <ENTRY entrytime="00:01:12.19" eventid="1785" heatid="4719" lane="2" />
                <ENTRY entrytime="00:01:12.21" eventid="1799" heatid="4732" lane="3" />
                <ENTRY entrytime="00:02:20.16" eventid="1978" heatid="4830" lane="2" />
                <ENTRY entrytime="00:00:33.91" eventid="2034" heatid="4884" lane="2" />
                <ENTRY entrytime="00:02:38.37" eventid="2055" heatid="4898" lane="1" />
                <ENTRY entrytime="00:02:33.79" eventid="2096" heatid="4933" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Gina" gender="F" lastname="Mayer" nation="GER" license="257249" athleteid="2721">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.02" eventid="1059" heatid="4670" lane="6" />
                <ENTRY entrytime="00:01:11.93" eventid="1799" heatid="4733" lane="4" />
                <ENTRY entrytime="00:04:48.88" eventid="1827" heatid="4761" lane="6" />
                <ENTRY entrytime="00:02:12.97" eventid="1978" heatid="4835" lane="1" />
                <ENTRY entrytime="00:00:32.66" eventid="2034" heatid="4886" lane="2" />
                <ENTRY entrytime="00:02:34.12" eventid="2055" heatid="4901" lane="6" />
                <ENTRY entrytime="00:00:28.84" eventid="2082" heatid="4918" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Wolfgang" gender="M" lastname="Orth" nation="GER" license="226633" athleteid="2729">
              <ENTRIES>
                <ENTRY entrytime="00:01:58.91" eventid="1749" heatid="4683" lane="6" />
                <ENTRY entrytime="00:16:27.61" eventid="1792" heatid="4727" lane="2" />
                <ENTRY entrytime="00:02:15.37" eventid="1848" heatid="4790" lane="6" />
                <ENTRY entrytime="00:00:55.62" eventid="1971" heatid="4821" lane="5" />
                <ENTRY entrytime="00:01:03.56" eventid="2013" heatid="4870" lane="2" />
                <ENTRY entrytime="00:04:11.03" eventid="2075" heatid="4911" lane="6" />
                <ENTRY entrytime="00:08:48.98" eventid="2168" heatid="4808" lane="6">
                  <MEETINFO qualificationtime="00:08:48.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Johannes" gender="M" lastname="Vorbach" nation="GER" license="257156" athleteid="2737">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.63" eventid="1763" heatid="4696" lane="3" />
                <ENTRY entrytime="00:00:27.37" eventid="1834" heatid="4765" lane="4" />
                <ENTRY entrytime="00:00:58.81" eventid="1971" heatid="4815" lane="6" />
                <ENTRY entrytime="00:00:33.61" eventid="1985" heatid="4842" lane="6" />
                <ENTRY entrytime="00:02:42.43" eventid="2089" heatid="4925" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Lea" gender="F" lastname="Wienstruck" nation="GER" license="296635" athleteid="2743">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.91" eventid="1059" heatid="4664" lane="4" />
                <ENTRY entrytime="00:01:10.27" eventid="1785" heatid="4721" lane="1" />
                <ENTRY entrytime="00:01:12.09" eventid="1799" heatid="4733" lane="1" />
                <ENTRY entrytime="00:00:32.59" eventid="2034" heatid="4886" lane="4" />
                <ENTRY entrytime="00:02:34.66" eventid="2055" heatid="4900" lane="3" />
                <ENTRY entrytime="00:00:29.22" eventid="2082" heatid="4916" lane="5" />
                <ENTRY entrytime="00:02:29.99" eventid="2096" heatid="4934" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4397" nation="GER" region="02" clubid="2751" name="TG Kitzingen">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Viktoria" gender="F" lastname="Kolb" nation="GER" license="291280" athleteid="2752">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.51" eventid="1059" heatid="4665" lane="3" />
                <ENTRY entrytime="00:01:14.51" eventid="1799" heatid="4729" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4405" nation="GER" region="02" clubid="4159" name="TSG Kleinostheim">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Francis" gender="M" lastname="Hartl" nation="GER" license="285486" athleteid="4163">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.09" eventid="1971" heatid="4813" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Alena" gender="F" lastname="Hennl" nation="GER" license="208754" athleteid="4165">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.93" eventid="1756" heatid="4693" lane="2" />
                <ENTRY entrytime="00:02:25.46" eventid="1813" heatid="4747" lane="2" />
                <ENTRY entrytime="00:00:29.91" eventid="1855" heatid="4801" lane="6" />
                <ENTRY entrytime="00:01:16.85" eventid="1992" heatid="4855" lane="6" />
                <ENTRY entrytime="00:01:05.46" eventid="2006" heatid="4866" lane="2" />
                <ENTRY entrytime="00:02:28.56" eventid="2055" heatid="4902" lane="1" />
                <ENTRY entrytime="00:00:33.58" eventid="1877" heatid="4695" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.26" eventid="1933" heatid="5429" lane="3">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.57" eventid="1940" heatid="5517" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4439" nation="GER" region="02" clubid="2481" name="TSV - Eintracht Karlsfeld">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Johannes" gender="M" lastname="Heizenreder" nation="GER" license="248442" athleteid="2482">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.25" eventid="1806" heatid="4741" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Miriam" gender="F" lastname="Zanklmaier" nation="GER" license="283818" athleteid="2484">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.50" eventid="1756" heatid="4690" lane="6" />
                <ENTRY entrytime="00:01:11.50" eventid="1799" heatid="4734" lane="1" />
                <ENTRY entrytime="00:00:30.50" eventid="1855" heatid="4799" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4413" nation="GER" region="02" clubid="2674" name="TSV 1860 Rosenheim">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Alexander" gender="M" lastname="Bauer" nation="GER" license="257560" athleteid="2675">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.58" eventid="1778" heatid="4711" lane="6" />
                <ENTRY entrytime="00:00:28.45" eventid="2103" heatid="4941" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Paula" gender="F" lastname="Borst" nation="GER" license="200640" athleteid="2678">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.90" eventid="1059" heatid="4670" lane="5" />
                <ENTRY entrytime="00:00:30.50" eventid="1855" heatid="4799" lane="4" />
                <ENTRY entrytime="00:00:28.20" eventid="2082" heatid="4922" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Lucas" gender="M" lastname="Kleinicke" nation="GER" license="226836" athleteid="2682">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.00" eventid="1749" heatid="4678" lane="1" />
                <ENTRY entrytime="00:01:01.20" eventid="1778" heatid="4712" lane="4" />
                <ENTRY entrytime="00:00:24.86" eventid="1834" heatid="4774" lane="5" />
                <ENTRY entrytime="00:00:57.20" eventid="1971" heatid="4818" lane="6" />
                <ENTRY entrytime="00:00:27.42" eventid="2103" heatid="4943" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Alexandra" gender="F" lastname="Schöne" nation="GER" license="266174" athleteid="2688">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.06" eventid="1059" heatid="4669" lane="3" />
                <ENTRY entrytime="00:01:08.87" eventid="1785" heatid="4721" lane="3" />
                <ENTRY entrytime="00:04:41.00" eventid="1827" heatid="4762" lane="5" />
                <ENTRY entrytime="00:02:12.25" eventid="1978" heatid="4835" lane="4" />
                <ENTRY entrytime="00:00:30.90" eventid="2034" heatid="4889" lane="2" />
                <ENTRY entrytime="00:00:28.30" eventid="2082" heatid="4920" lane="2" />
                <ENTRY entrytime="00:02:33.62" eventid="2096" heatid="4933" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Sarah" gender="F" lastname="Wieser" nation="GER" license="295252" athleteid="2696">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.07" eventid="1855" heatid="4794" lane="5" />
                <ENTRY entrytime="00:00:34.27" eventid="2034" heatid="4883" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4441" nation="GER" region="02" clubid="3253" name="TSV Erding">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Carina" gender="F" lastname="Michaelis" nation="GER" license="313153" athleteid="3254">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.17" eventid="1059" heatid="4666" lane="3" />
                <ENTRY entrytime="00:01:12.64" eventid="1799" heatid="4732" lane="6" />
                <ENTRY entrytime="00:04:55.07" eventid="1827" heatid="4758" lane="3" />
                <ENTRY entrytime="00:00:30.67" eventid="1855" heatid="4799" lane="1" />
                <ENTRY entrytime="00:02:15.65" eventid="1978" heatid="4833" lane="5" />
                <ENTRY entrytime="00:00:33.97" eventid="2034" heatid="4884" lane="5" />
                <ENTRY entrytime="00:02:37.06" eventid="2055" heatid="4899" lane="1" />
                <ENTRY entrytime="00:00:28.97" eventid="2082" heatid="4917" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4452" nation="GER" region="02" clubid="2771" name="TSV Hohenbrunn-Riemerl.">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Nick" gender="M" lastname="Bongartz" nation="GER" license="325785" athleteid="2772">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.58" eventid="1749" heatid="4679" lane="5" />
                <ENTRY entrytime="00:02:20.68" eventid="1820" heatid="4752" lane="1" />
                <ENTRY entrytime="00:00:57.45" eventid="1971" heatid="4817" lane="4" />
                <ENTRY entrytime="00:05:02.54" eventid="1999" heatid="4860" lane="2" />
                <ENTRY entrytime="00:04:33.74" eventid="2075" heatid="4908" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Adrien" gender="M" lastname="Cara" nation="GER" license="294598" athleteid="2778">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.44" eventid="1763" heatid="4697" lane="5" />
                <ENTRY entrytime="00:02:22.77" eventid="1820" heatid="4750" lane="3" />
                <ENTRY entrytime="00:02:17.35" eventid="1848" heatid="4788" lane="3" />
                <ENTRY entrytime="00:00:57.50" eventid="1971" heatid="4817" lane="2" />
                <ENTRY entrytime="00:04:59.19" eventid="1999" heatid="4860" lane="4" />
                <ENTRY entrytime="00:01:03.36" eventid="2013" heatid="4870" lane="3" />
                <ENTRY entrytime="00:02:38.40" eventid="2089" heatid="4926" lane="5" />
                <ENTRY entrytime="00:02:16.91" eventid="1961" heatid="5504" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Daniela" gender="F" lastname="Ernst" nation="GER" license="316890" athleteid="2786">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.57" eventid="1785" heatid="4720" lane="1" />
                <ENTRY entrytime="00:00:33.98" eventid="2034" heatid="4884" lane="1" />
                <ENTRY entrytime="00:02:32.23" eventid="2096" heatid="4934" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lisa-Marie" gender="F" lastname="Geisler" nation="GER" license="221272" athleteid="2790">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.03" eventid="1756" heatid="4690" lane="4" />
                <ENTRY entrytime="00:02:49.25" eventid="1841" heatid="4781" lane="4" />
                <ENTRY entrytime="00:01:17.28" eventid="1992" heatid="4854" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Amna" gender="F" lastname="Hasanbegovic" nation="GER" license="225371" athleteid="2794">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.80" eventid="1799" heatid="4731" lane="4" />
                <ENTRY entrytime="00:00:31.08" eventid="1855" heatid="4797" lane="1" />
                <ENTRY entrytime="00:01:08.34" eventid="2006" heatid="4865" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Eric Florian" gender="M" lastname="Henschel" nation="GER" license="212691" athleteid="2798">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.66" eventid="1834" heatid="4771" lane="1" />
                <ENTRY entrytime="00:00:56.98" eventid="1971" heatid="4818" lane="5" />
                <ENTRY entrytime="00:00:27.42" eventid="2103" heatid="4943" lane="3" />
                <ENTRY entrytime="00:00:24.23" eventid="1947" heatid="5478" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Alina" gender="F" lastname="Hermeking" nation="GER" license="290265" athleteid="2802">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.33" eventid="1756" heatid="4688" lane="2" />
                <ENTRY entrytime="00:01:22.48" eventid="1992" heatid="4850" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Fabian" gender="M" lastname="Hoffmann" nation="GER" license="290269" athleteid="2805">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.05" eventid="1806" heatid="4738" lane="3" />
                <ENTRY entrytime="00:00:26.46" eventid="1834" heatid="4768" lane="1" />
                <ENTRY entrytime="00:00:59.46" eventid="1971" heatid="4814" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Tobias" gender="M" lastname="Hollaus" nation="GER" license="209181" athleteid="2809">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.32" eventid="1763" heatid="4702" lane="2" />
                <ENTRY entrytime="00:00:29.90" eventid="1985" heatid="4848" lane="5" />
                <ENTRY entrytime="00:02:22.45" eventid="2089" heatid="4928" lane="4" />
                <ENTRY entrytime="00:01:04.10" eventid="1884" heatid="4704" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Sarah-Isabelle" gender="F" lastname="Mai" nation="GER" license="269795" athleteid="2813">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.56" eventid="1756" heatid="4693" lane="5" />
                <ENTRY entrytime="00:01:09.56" eventid="1799" heatid="4736" lane="5" />
                <ENTRY entrytime="00:02:45.89" eventid="1841" heatid="4783" lane="1" />
                <ENTRY entrytime="00:01:15.81" eventid="1992" heatid="4856" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1994-01-01" firstname="Francesco" gender="M" lastname="Montanari" nation="GER" license="281775" athleteid="2818">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.94" eventid="1834" heatid="4773" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Tom" gender="M" lastname="Nolte" nation="GER" license="288931" athleteid="2820">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.77" eventid="1763" heatid="4698" lane="6" />
                <ENTRY entrytime="00:00:30.16" eventid="1806" heatid="4739" lane="3" />
                <ENTRY entrytime="00:00:25.92" eventid="1834" heatid="4770" lane="2" />
                <ENTRY entrytime="00:00:32.81" eventid="1985" heatid="4842" lane="2" />
                <ENTRY entrytime="00:01:06.15" eventid="2013" heatid="4869" lane="2" />
                <ENTRY entrytime="00:00:28.85" eventid="2103" heatid="4940" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Sven" gender="M" lastname="Pesut" nation="GER" license="360757" athleteid="2827">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.16" eventid="1749" heatid="4680" lane="6" />
                <ENTRY entrytime="00:01:01.85" eventid="1778" heatid="4712" lane="6" />
                <ENTRY entrytime="00:02:22.35" eventid="1820" heatid="4751" lane="1" />
                <ENTRY entrytime="00:00:56.72" eventid="1971" heatid="4819" lane="3" />
                <ENTRY entrytime="00:05:06.39" eventid="1999" heatid="4859" lane="4" />
                <ENTRY entrytime="00:04:31.63" eventid="2075" heatid="4908" lane="2" />
                <ENTRY entrytime="00:00:27.56" eventid="2103" heatid="4943" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Noah" gender="M" lastname="Rueff" nation="GER" license="241485" athleteid="2835">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.80" eventid="1778" heatid="4710" lane="3" />
                <ENTRY entrytime="00:00:30.30" eventid="1806" heatid="4739" lane="2" />
                <ENTRY entrytime="00:00:33.00" eventid="1985" heatid="4842" lane="5" />
                <ENTRY entrytime="00:01:05.20" eventid="2013" heatid="4869" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Moritz" gender="M" lastname="Schepp" nation="GER" license="279390" athleteid="2840">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.27" eventid="1806" heatid="4739" lane="4" />
                <ENTRY entrytime="00:00:26.33" eventid="1834" heatid="4768" lane="2" />
                <ENTRY entrytime="00:02:20.87" eventid="1848" heatid="4787" lane="4" />
                <ENTRY entrytime="00:00:58.07" eventid="1971" heatid="4816" lane="1" />
                <ENTRY entrytime="00:01:06.39" eventid="2013" heatid="4869" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Florian" gender="M" lastname="Schimanski" nation="GER" license="183469" athleteid="2846">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.64" eventid="1778" heatid="4713" lane="4" />
                <ENTRY entrytime="00:00:24.94" eventid="1834" heatid="4774" lane="6" />
                <ENTRY entrytime="00:00:54.07" eventid="1971" heatid="4824" lane="2" />
                <ENTRY entrytime="00:00:25.60" eventid="2103" heatid="4947" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Nico" gender="M" lastname="Schmid" nation="GER" license="175732" athleteid="2851">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.23" eventid="1749" heatid="4685" lane="6" />
                <ENTRY entrytime="00:02:09.60" eventid="1820" heatid="4755" lane="2" />
                <ENTRY entrytime="00:00:24.63" eventid="1834" heatid="4775" lane="6" />
                <ENTRY entrytime="00:04:35.89" eventid="1999" heatid="4862" lane="2" />
                <ENTRY entrytime="00:04:08.23" eventid="2075" heatid="4911" lane="4" />
                <ENTRY entrytime="NT" eventid="2168" status="RJC" />
                <ENTRY entrytime="00:01:57.24" eventid="1870" heatid="5342" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.29" eventid="1926" heatid="5442" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Magnus" gender="M" lastname="Schweiger" nation="GER" license="158545" athleteid="2858">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.87" eventid="1749" heatid="4685" lane="2" />
                <ENTRY entrytime="00:00:58.90" eventid="1778" heatid="4716" lane="5" />
                <ENTRY entrytime="00:00:53.55" eventid="1971" heatid="4826" lane="6" />
                <ENTRY entrytime="00:02:10.69" eventid="2041" heatid="4893" lane="2" />
                <ENTRY entrytime="00:04:03.77" eventid="2075" heatid="4912" lane="6" />
                <ENTRY entrytime="00:01:54.03" eventid="1870" heatid="4686" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.93" eventid="1898" heatid="4717" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Helena" gender="F" lastname="Sedlar" nation="GER" license="290267" athleteid="2864">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.91" eventid="1059" heatid="4667" lane="5" />
                <ENTRY entrytime="00:04:55.05" eventid="1827" heatid="4759" lane="1" />
                <ENTRY entrytime="00:00:31.78" eventid="1855" heatid="4795" lane="1" />
                <ENTRY entrytime="00:02:21.10" eventid="1978" heatid="4829" lane="2" />
                <ENTRY entrytime="00:00:30.03" eventid="2082" heatid="4913" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lana" gender="F" lastname="Sokac" nation="GER" license="360313" athleteid="2870">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.83" eventid="1059" heatid="4674" lane="2" />
                <ENTRY entrytime="00:01:07.60" eventid="1799" heatid="4736" lane="2" />
                <ENTRY entrytime="00:00:29.35" eventid="1855" heatid="4801" lane="2" />
                <ENTRY entrytime="00:01:06.20" eventid="2006" heatid="4867" lane="5" />
                <ENTRY entrytime="00:00:26.68" eventid="2082" heatid="4922" lane="3" />
                <ENTRY entrytime="00:00:58.97" eventid="1863" heatid="4675" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.42" eventid="1919" heatid="4737" lane="1">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.92" eventid="1940" heatid="4802" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Jacopo" gender="M" lastname="Vercelli" nation="GER" license="329282" athleteid="2876">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.59" eventid="1778" heatid="4709" lane="5" />
                <ENTRY entrytime="00:00:26.70" eventid="1834" heatid="4767" lane="4" />
                <ENTRY entrytime="00:00:58.50" eventid="1971" heatid="4815" lane="5" />
                <ENTRY entrytime="00:02:24.00" eventid="2041" heatid="4891" lane="2" />
                <ENTRY entrytime="00:00:29.00" eventid="2103" heatid="4939" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Sina" gender="F" lastname="Wappenschmidt" nation="GER" license="269801" swrid="4642730" athleteid="2882">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.74" eventid="1059" heatid="4667" lane="3" />
                <ENTRY entrytime="00:01:10.96" eventid="1785" heatid="4720" lane="4" />
                <ENTRY entrytime="00:04:46.45" eventid="1827" heatid="4761" lane="5" />
                <ENTRY entrytime="00:19:00.94" eventid="1905" status="RJC">
                  <MEETINFO qualificationtime="00:19:00.94" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.63" eventid="1978" heatid="4832" lane="1" />
                <ENTRY entrytime="00:02:33.79" eventid="2055" heatid="4901" lane="2" />
                <ENTRY entrytime="00:02:33.74" eventid="2096" heatid="4933" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Florian" gender="M" lastname="Wutz" nation="GER" license="233903" athleteid="2890">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.16" eventid="1749" heatid="4681" lane="2" />
                <ENTRY entrytime="00:00:26.17" eventid="1834" heatid="4769" lane="5" />
                <ENTRY entrytime="00:00:57.34" eventid="1971" heatid="4817" lane="3" />
                <ENTRY entrytime="00:04:22.04" eventid="2075" heatid="4909" lane="4" />
                <ENTRY entrytime="00:09:20.58" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:20.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Niklas" gender="M" lastname="Zimmermann" nation="GER" license="345171" athleteid="2896">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.95" eventid="1763" heatid="4700" lane="5" />
                <ENTRY entrytime="00:00:26.26" eventid="1834" heatid="4769" lane="1" />
                <ENTRY entrytime="00:00:31.68" eventid="1985" heatid="4844" lane="4" />
                <ENTRY entrytime="00:02:31.33" eventid="2089" heatid="4927" lane="4" />
                <ENTRY entrytime="00:00:28.55" eventid="2103" heatid="4941" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.00" eventid="2048" heatid="4806" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2851" number="1" />
                    <RELAYPOSITION athleteid="2809" number="2" />
                    <RELAYPOSITION athleteid="2846" number="3" />
                    <RELAYPOSITION athleteid="2798" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:40.00" eventid="2232" heatid="4812" lane="1" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="2062" heatid="4807" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2786" number="1" />
                    <RELAYPOSITION athleteid="2813" number="2" />
                    <RELAYPOSITION athleteid="2794" number="3" />
                    <RELAYPOSITION athleteid="2870" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:55.00" eventid="2224" heatid="4810" lane="5" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4420" nation="GER" region="02" clubid="3434" name="TSV Neuburg">
          <ATHLETES>
            <ATHLETE birthdate="1979-01-01" firstname="Fabian" gender="M" lastname="Rieß" nation="GER" license="363828" athleteid="3440">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.97" eventid="1778" heatid="4714" lane="1" />
                <ENTRY entrytime="00:00:27.60" eventid="1806" heatid="4741" lane="4" />
                <ENTRY entrytime="00:02:15.14" eventid="1848" heatid="4789" lane="1" />
                <ENTRY entrytime="00:00:54.19" eventid="1971" heatid="4824" lane="1" />
                <ENTRY entrytime="00:01:00.26" eventid="2013" heatid="4873" lane="2" />
                <ENTRY entrytime="00:00:26.43" eventid="2103" heatid="4945" lane="5" />
                <ENTRY entrytime="00:00:27.22" eventid="1912" heatid="4744" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.90" eventid="1898" heatid="5465" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Christina" gender="F" lastname="Wenger" nation="GER" license="162995" athleteid="3435">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.77" eventid="1756" heatid="4692" lane="1" />
                <ENTRY entrytime="00:01:12.08" eventid="1799" heatid="4733" lane="5" />
                <ENTRY entrytime="00:00:31.05" eventid="1855" heatid="4797" lane="5" />
                <ENTRY entrytime="00:01:16.16" eventid="1992" heatid="4855" lane="5" />
                <ENTRY entrytime="00:00:34.66" eventid="1877" heatid="5355" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4492" nation="GER" region="02" clubid="3786" name="TSV Vaterstetten">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Christian" gender="M" lastname="Arzberger" nation="GER" license="290446" athleteid="3785">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.80" eventid="1985" heatid="4840" lane="2" />
                <ENTRY entrytime="00:02:42.51" eventid="2089" heatid="4925" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Pauline" gender="F" lastname="Breitner" nation="GER" license="273792" athleteid="3789">
              <ENTRIES>
                <ENTRY entrytime="00:02:20.01" eventid="1978" heatid="4830" lane="4" />
                <ENTRY entrytime="00:01:20.60" eventid="1992" heatid="4851" lane="5" />
                <ENTRY entrytime="00:02:40.29" eventid="2055" heatid="4896" lane="1" />
                <ENTRY entrytime="00:00:29.54" eventid="2082" heatid="4914" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Valerie" gender="F" lastname="Wende" nation="GER" license="325391" athleteid="3794">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.65" eventid="2082" heatid="4914" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5107" nation="GER" region="02" clubid="2650" name="TV 1860 Immenstadt">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Marcus" gender="M" lastname="Joas" nation="GER" license="161806" athleteid="2651">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1749" heatid="4679" lane="2" />
                <ENTRY entrytime="00:02:22.29" eventid="1820" heatid="4751" lane="5" />
                <ENTRY entrytime="00:02:21.68" eventid="1848" heatid="4787" lane="1" />
                <ENTRY entrytime="00:00:58.10" eventid="1971" heatid="4815" lane="4" />
                <ENTRY entrytime="00:02:21.10" eventid="2041" heatid="4891" lane="4" />
                <ENTRY entrytime="00:04:22.25" eventid="2075" heatid="4909" lane="5" />
                <ENTRY entrytime="00:08:58.39" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:08:58.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Simon" gender="M" lastname="Joas" nation="GER" license="282570" athleteid="2659">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.06" eventid="1749" heatid="4677" lane="2" />
                <ENTRY entrytime="00:00:27.34" eventid="1834" heatid="4766" lane="5" />
                <ENTRY entrytime="00:00:59.59" eventid="1971" heatid="4814" lane="5" />
                <ENTRY entrytime="00:04:34.09" eventid="2075" heatid="4907" lane="3" />
                <ENTRY entrytime="00:09:23.29" eventid="2168" status="RJC">
                  <MEETINFO qualificationtime="00:09:23.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4530" nation="GER" region="02" clubid="2495" name="TV 1862 Passau">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Luisa" gender="F" lastname="Roderweis" nation="GER" license="245436" athleteid="2496">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.57" eventid="1785" heatid="4724" lane="1" />
                <ENTRY entrytime="00:02:23.87" eventid="1813" heatid="4745" lane="4" />
                <ENTRY entrytime="00:04:25.65" eventid="1827" heatid="4764" lane="5" />
                <ENTRY entrytime="00:02:07.47" eventid="1978" heatid="4838" lane="2" />
                <ENTRY entrytime="00:09:19.00" eventid="2020" heatid="4876" lane="5">
                  <MEETINFO qualificationtime="00:09:18.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.32" eventid="2096" heatid="4936" lane="2" />
                <ENTRY entrytime="00:01:06.65" eventid="1891" heatid="5391" lane="5">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.69" eventid="1933" heatid="4748" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6812" nation="GER" region="02" clubid="2411" name="TV Kempten">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Jannes" gender="M" lastname="Schnitzer" nation="GER" license="294908" athleteid="2412">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.94" eventid="1763" heatid="4700" lane="6" />
                <ENTRY entrytime="00:01:00.96" eventid="1778" heatid="4713" lane="5" />
                <ENTRY entrytime="00:02:16.61" eventid="1820" heatid="4753" lane="6" />
                <ENTRY entrytime="00:02:18.28" eventid="1848" heatid="4788" lane="2" />
                <ENTRY entrytime="00:00:32.53" eventid="1985" heatid="4843" lane="1" />
                <ENTRY entrytime="00:01:00.67" eventid="2013" heatid="4872" lane="2" />
                <ENTRY entrytime="00:01:03.52" eventid="2027" heatid="4879" lane="6" />
                <ENTRY entrytime="00:02:18.14" eventid="2041" heatid="4893" lane="6" />
                <ENTRY entrytime="00:02:36.99" eventid="2089" heatid="4926" lane="4" />
                <ENTRY entrytime="00:02:15.55" eventid="1961" heatid="5504" lane="4">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Jan" gender="M" lastname="Schuster" nation="GER" license="301516" athleteid="2422">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.14" eventid="1749" heatid="4678" lane="2" />
                <ENTRY entrytime="00:01:02.20" eventid="1778" heatid="4711" lane="5" />
                <ENTRY entrytime="00:00:30.31" eventid="1806" heatid="4739" lane="5" />
                <ENTRY entrytime="00:00:25.78" eventid="1834" heatid="4770" lane="3" />
                <ENTRY entrytime="00:00:56.68" eventid="1971" heatid="4820" lane="6" />
                <ENTRY entrytime="00:01:05.05" eventid="2027" heatid="4878" lane="5" />
                <ENTRY entrytime="00:00:27.07" eventid="2103" heatid="4944" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Lucas" gender="M" lastname="Willinsky" nation="GER" license="248935" athleteid="2430">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.50" eventid="1763" heatid="4701" lane="2" />
                <ENTRY entrytime="00:00:28.96" eventid="1806" heatid="4741" lane="1" />
                <ENTRY entrytime="00:00:29.80" eventid="1985" heatid="4846" lane="2" />
                <ENTRY entrytime="00:01:01.14" eventid="2027" heatid="4879" lane="2" />
                <ENTRY entrytime="00:02:21.88" eventid="2089" heatid="4929" lane="4" />
                <ENTRY entrytime="00:01:04.52" eventid="1884" heatid="5368" lane="2">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.69" eventid="1912" heatid="5417" lane="6">
                  <MEETINFO qualificationtime="00:00:00.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4562" nation="GER" region="02" clubid="3230" name="TV Parsberg">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Alicia" gender="F" lastname="Urschel" nation="GER" license="300240" athleteid="3231">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.08" eventid="1059" heatid="4669" lane="4" />
                <ENTRY entrytime="00:05:40.46" eventid="1771" heatid="4705" lane="2" />
                <ENTRY entrytime="00:01:13.63" eventid="1799" heatid="4730" lane="1" />
                <ENTRY entrytime="00:02:18.47" eventid="1978" heatid="4831" lane="3" />
                <ENTRY entrytime="00:02:39.55" eventid="2055" heatid="4896" lane="4" />
                <ENTRY entrytime="00:00:28.43" eventid="2082" heatid="4919" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4593" nation="GER" region="02" clubid="4270" name="VfL 1860 Spfr. Bad Neustadt">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Sebastian" gender="M" lastname="Rasch" nation="GER" license="305639" athleteid="4569">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.45" eventid="1834" heatid="4768" lane="5" />
                <ENTRY entrytime="00:00:57.94" eventid="1971" heatid="4816" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1062" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="15" agemin="-1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:25.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:24.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:43.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.20">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:28.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:16.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:16.90">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1064" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="15" agemin="-1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:38.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:37.60">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:58.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:21.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:59.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:14.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.90">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:41.50">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1066" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:25.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:24.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:43.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:40.20">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:07.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:28.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:16.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:16.90">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1068" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:37.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.20">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:56.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:55.20">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:39.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:21.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:38.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:14.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1078" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="18" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:22.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:21.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:38.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:07.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:31.70">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:23.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:09.10">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1080" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="18" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:32.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:32.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:51.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:49.70">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:19.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:31.80">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1070" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="19" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:18.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:33.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:04.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:25.10">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:01.80">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:01.40">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:04.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1072" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="19" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:32.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:32.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:51.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:49.70">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:19.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:31.80">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="2070" code="BAY" course="SCM" gender="M" name="Bayerische Kurzbahn Staffel" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:47.50">
          <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:15.00">
          <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="2072" code="BAY" course="SCM" gender="F" name="Bayerische Kurzbahn Staffel" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
