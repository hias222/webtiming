<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SG Fürth" version="11.61084">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Nürnberg" name="Bayerische Kurzbahnmeisterschaften 2019" course="SCM" deadline="2019-10-14" hostclub="TSV Altenfurt Nürnberg" organizer="Bayerischer Schwimmverband" organizer.url="https://www.bayerischer-schwimmverband.de" reservecount="6" startmethod="1" timing="AUTOMATIC" withdrawuntil="2019-10-16" nation="GER">
      <AGEDATE value="2019-10-20" type="YEAR" />
      <POOL name="Hallenbad Langwasser" lanemin="1" lanemax="6" />
      <FACILITY city="Nürnberg" name="Hallenbad Langwasser" nation="GER" street="Breslauer Straße 251" zip="90471" />
      <POINTTABLE pointtableid="3012" name="FINA Point Scoring" version="2019" />
      <CONTACT email="meldungen@sgfuerth.de" name="Matthias Fuchs" phone="09118101172" />
      <QUALIFY from="2019-01-01" until="2019-10-18" conversion="NON_CONFORMING_LAST" />
      <SESSIONS>
        <SESSION date="2019-10-19" daytime="10:00" number="1" officialmeeting="09:00" teamleadermeeting="09:00" warmupfrom="08:30" warmupuntil="09:50">
          <EVENTS>
            <EVENT eventid="1841" daytime="13:25" gender="F" number="15" order="15" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9457" daytime="13:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9458" daytime="13:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9459" daytime="13:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9460" daytime="13:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9461" daytime="13:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9462" daytime="13:30" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9463" daytime="13:30" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1059" daytime="10:00" gender="F" number="1" order="1" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9345" daytime="10:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9346" daytime="10:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9347" daytime="10:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9348" daytime="10:05" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9349" daytime="10:05" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9350" daytime="10:10" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9351" daytime="10:10" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9352" daytime="10:10" number="8" order="8" status="SEEDED" />
                <HEAT heatid="9353" daytime="10:10" number="9" order="9" status="SEEDED" />
                <HEAT heatid="9354" daytime="10:15" number="10" order="10" status="SEEDED" />
                <HEAT heatid="9355" daytime="10:15" number="11" order="11" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1763" daytime="10:45" gender="M" number="4" order="4" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9377" daytime="10:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9378" daytime="10:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9379" daytime="10:50" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9380" daytime="10:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9381" daytime="10:55" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9382" daytime="10:55" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9383" daytime="10:55" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9384" daytime="11:00" number="8" order="8" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1813" daytime="12:35" gender="F" number="11" order="11" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9425" daytime="12:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9426" daytime="12:40" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1848" daytime="13:30" gender="M" number="16" order="16" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9466" daytime="13:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9467" daytime="13:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9468" daytime="13:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9469" daytime="13:40" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1771" daytime="11:00" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9387" daytime="11:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9388" daytime="11:05" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1792" daytime="11:35" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9406" daytime="11:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9407" daytime="12:00" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1855" daytime="14:05" gender="X" number="18" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="2500" />
              <HEATS>
                <HEAT heatid="9476" daytime="14:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9477" daytime="14:10" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1827" daytime="13:00" gender="F" number="13" order="13" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9436" daytime="13:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9437" daytime="13:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9438" daytime="13:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9439" daytime="13:10" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1799" daytime="12:15" gender="F" number="9" order="9" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9408" daytime="12:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9409" daytime="12:20" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9410" daytime="12:20" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9411" daytime="12:20" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9412" daytime="12:25" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9413" daytime="12:25" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9414" daytime="12:25" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9415" daytime="12:30" number="8" order="8" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1820" daytime="12:45" gender="M" number="12" order="12" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9429" daytime="12:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9430" daytime="12:45" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9431" daytime="12:50" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9432" daytime="12:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9433" daytime="12:55" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1756" daytime="10:40" gender="F" number="3" order="3" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9368" daytime="10:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9369" daytime="10:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9370" daytime="10:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9371" daytime="10:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9372" daytime="10:45" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9373" daytime="10:45" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9374" daytime="10:45" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1834" daytime="13:10" gender="M" number="14" order="14" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9442" daytime="13:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9443" daytime="13:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9444" daytime="13:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9445" daytime="13:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9446" daytime="13:15" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9447" daytime="13:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9448" daytime="13:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9449" daytime="13:20" number="8" order="8" status="SEEDED" />
                <HEAT heatid="9450" daytime="13:20" number="9" order="9" status="SEEDED" />
                <HEAT heatid="9451" daytime="13:20" number="10" order="10" status="SEEDED" />
                <HEAT heatid="9452" daytime="13:20" number="11" order="11" status="SEEDED" />
                <HEAT heatid="9453" daytime="13:20" number="12" order="12" status="SEEDED" />
                <HEAT heatid="9454" daytime="13:25" number="13" order="13" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1785" daytime="11:25" gender="F" number="7" order="7" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9397" daytime="11:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9398" daytime="11:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9399" daytime="11:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9400" daytime="11:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9401" daytime="11:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9402" daytime="11:30" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9403" daytime="11:35" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1749" daytime="10:15" gender="M" number="2" order="2" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9358" daytime="10:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9359" daytime="10:20" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9360" daytime="10:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9361" daytime="10:25" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9362" daytime="10:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9363" daytime="10:30" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9364" daytime="10:35" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9365" daytime="10:35" number="8" order="8" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5320" daytime="13:45" gender="F" number="17" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9472" daytime="13:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9473" daytime="13:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9474" daytime="13:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9475" daytime="14:00" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1806" daytime="12:30" gender="M" number="10" order="10" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9418" daytime="12:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9419" daytime="12:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9420" daytime="12:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9421" daytime="12:35" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9422" daytime="12:35" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1778" daytime="11:15" gender="M" number="6" order="6" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9389" daytime="11:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9390" daytime="11:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9391" daytime="11:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9392" daytime="11:20" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9393" daytime="11:20" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9394" daytime="11:20" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-10-19" daytime="16:00" number="2">
          <EVENTS>
            <EVENT eventid="7586" gender="M" number="10" order="8" round="FIN" preveventid="1806">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="9423" agegroupid="7587" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9424" agegroupid="7587" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7596" gender="M" number="12" order="10" round="FIN" preveventid="1820">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="9434" agegroupid="7597" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9435" agegroupid="7597" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5314" gender="F" number="21" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="2500" />
              <HEATS>
                <HEAT heatid="9482" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9483" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7616" gender="M" number="16" order="14" round="FIN" preveventid="1848">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="9470" agegroupid="7617" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9471" agegroupid="7617" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5318" gender="F" number="19" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9478" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9479" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7601" gender="F" number="13" order="13" round="FIN" preveventid="1827">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="9440" agegroupid="7602" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9441" agegroupid="7602" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7551" gender="M" number="2" order="2" round="FIN" preveventid="1749">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="9366" agegroupid="7552" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9367" agegroupid="7552" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7576" gender="F" number="7" order="5" round="FIN" preveventid="1785">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="9404" agegroupid="7577" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9405" agegroupid="7577" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5316" gender="M" number="20" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="2500" />
              <HEATS>
                <HEAT heatid="9480" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9481" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7556" gender="F" number="3" order="3" round="FIN" preveventid="1756">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="9375" agegroupid="7557" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9376" agegroupid="7557" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7606" gender="M" number="14" order="12" round="FIN" preveventid="1834">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="9455" agegroupid="7607" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9456" agegroupid="7607" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7571" gender="M" number="6" order="6" round="FIN" preveventid="1778">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="9395" agegroupid="7572" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9396" agegroupid="7572" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7591" gender="F" number="11" order="11" round="FIN" preveventid="1813">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="9427" agegroupid="7592" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9428" agegroupid="7592" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7561" gender="M" number="4" order="4" round="FIN" preveventid="1763">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="9385" agegroupid="7562" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9386" agegroupid="7562" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5809" gender="F" number="1" order="1" round="FIN" preveventid="1059">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="9356" agegroupid="5810" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9357" agegroupid="5810" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7581" gender="F" number="9" order="9" round="FIN" preveventid="1799">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="9416" agegroupid="7582" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9417" agegroupid="7582" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7611" gender="F" number="15" order="15" round="FIN" preveventid="1841">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="9464" agegroupid="7612" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9465" agegroupid="7612" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-10-20" daytime="09:30" number="3" officialmeeting="09:00" teamleadermeeting="09:00" warmupfrom="07:45" warmupuntil="09:15">
          <EVENTS>
            <EVENT eventid="1999" daytime="10:30" gender="M" number="26" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9527" daytime="10:30" number="1" order="1" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2006" daytime="10:35" gender="F" number="27" order="6" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9528" daytime="10:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9529" daytime="10:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9530" daytime="10:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9531" daytime="10:40" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2041" daytime="11:20" gender="M" number="32" order="11" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9558" daytime="11:20" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9559" daytime="11:25" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2082" daytime="11:45" gender="M" number="34" order="13" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9570" daytime="11:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9571" daytime="11:50" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9572" daytime="11:50" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9573" daytime="11:55" number="4" order="4" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5307" daytime="12:10" gender="M" number="36" order="15" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9591" daytime="12:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9592" daytime="12:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9593" daytime="12:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9594" daytime="12:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9595" daytime="12:15" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9596" daytime="12:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9597" daytime="12:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9598" daytime="12:20" number="8" order="8" status="SEEDED" />
                <HEAT heatid="9599" daytime="12:20" number="9" order="9" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1971" daytime="09:30" gender="M" number="22" order="1" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9484" daytime="09:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9485" daytime="09:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9486" daytime="09:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9487" daytime="09:35" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9488" daytime="09:35" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9489" daytime="09:35" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9490" daytime="09:40" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9491" daytime="09:40" number="8" order="8" status="SEEDED" />
                <HEAT heatid="9492" daytime="09:40" number="9" order="9" status="SEEDED" />
                <HEAT heatid="9493" daytime="09:45" number="10" order="10" status="SEEDED" />
                <HEAT heatid="9494" daytime="09:45" number="11" order="11" status="SEEDED" />
                <HEAT heatid="9495" daytime="09:45" number="12" order="12" status="SEEDED" />
                <HEAT heatid="9496" daytime="09:45" number="13" order="13" status="SEEDED" />
                <HEAT heatid="9497" daytime="09:50" number="14" order="14" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2096" daytime="12:20" gender="F" number="37" order="16" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9602" daytime="12:20" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9603" daytime="12:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9604" daytime="12:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9605" daytime="12:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9606" daytime="12:35" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1985" daytime="10:10" gender="M" number="24" order="3" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9509" daytime="10:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9510" daytime="10:10" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9511" daytime="10:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9512" daytime="10:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9513" daytime="10:15" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9514" daytime="10:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9515" daytime="10:15" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9516" daytime="10:20" number="8" order="8" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2027" daytime="11:05" gender="M" number="30" order="9" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9542" daytime="11:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9543" daytime="11:05" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9544" daytime="11:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9545" daytime="11:10" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9546" daytime="11:10" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2013" daytime="10:45" gender="M" number="28" order="7" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9534" daytime="10:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9535" daytime="10:45" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9536" daytime="10:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9537" daytime="10:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9538" daytime="10:50" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2089" daytime="12:00" gender="F" number="35" order="14" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9576" daytime="12:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9577" daytime="12:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9578" daytime="12:00" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9579" daytime="12:00" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9580" daytime="12:00" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9581" daytime="12:05" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9582" daytime="12:05" number="7" order="7" status="SEEDED" />
                <HEAT heatid="9583" daytime="12:05" number="8" order="8" status="SEEDED" />
                <HEAT heatid="9584" daytime="12:05" number="9" order="9" status="SEEDED" />
                <HEAT heatid="9585" daytime="12:05" number="10" order="10" status="SEEDED" />
                <HEAT heatid="9586" daytime="12:10" number="11" order="11" status="SEEDED" />
                <HEAT heatid="9587" daytime="12:10" number="12" order="12" status="SEEDED" />
                <HEAT heatid="9588" daytime="12:10" number="13" order="13" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1978" daytime="09:50" gender="F" number="23" order="2" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9500" daytime="09:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9501" daytime="09:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9502" daytime="09:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9503" daytime="10:00" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9504" daytime="10:00" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9505" daytime="10:05" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9506" daytime="10:10" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1992" daytime="10:20" gender="F" number="25" order="4" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9519" daytime="10:20" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9520" daytime="10:20" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9521" daytime="10:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9522" daytime="10:25" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9523" daytime="10:25" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9524" daytime="10:30" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2020" daytime="10:50" gender="F" number="29" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9541" daytime="10:50" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2075" daytime="11:25" gender="F" number="33" order="12" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9562" daytime="11:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9563" daytime="11:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9564" daytime="11:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9565" daytime="11:35" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9566" daytime="11:40" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9567" daytime="11:40" number="6" order="6" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="5303" daytime="13:00" gender="X" number="39" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="2500" />
              <HEATS>
                <HEAT heatid="9614" daytime="13:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9615" daytime="13:05" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2034" daytime="11:10" gender="F" number="31" order="10" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9549" daytime="11:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9550" daytime="11:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9551" daytime="11:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9552" daytime="11:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9553" daytime="11:15" number="5" order="5" status="SEEDED" />
                <HEAT heatid="9554" daytime="11:20" number="6" order="6" status="SEEDED" />
                <HEAT heatid="9555" daytime="11:20" number="7" order="7" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2103" daytime="12:35" gender="M" number="38" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9609" daytime="12:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9610" daytime="12:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="9611" daytime="12:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="9612" daytime="12:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="9613" daytime="12:55" number="5" order="5" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-10-20" daytime="14:30" number="4">
          <EVENTS>
            <EVENT eventid="7646" gender="M" number="28" order="5" round="FIN" preveventid="2013">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="9539" agegroupid="7647" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9540" agegroupid="7647" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7621" gender="M" number="22" order="1" round="FIN" preveventid="1971">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="9498" agegroupid="7622" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9499" agegroupid="7622" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7661" gender="M" number="32" order="11" round="FIN" preveventid="2041">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="9560" agegroupid="7662" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9561" agegroupid="7662" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2168" gender="M" number="40" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="1200" />
              <HEATS>
                <HEAT heatid="9616" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9617" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7636" gender="F" number="25" order="4" round="FIN" preveventid="1992">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="9525" agegroupid="7637" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9526" agegroupid="7637" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7686" gender="F" number="37" order="14" round="FIN" preveventid="2096">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="9607" agegroupid="7687" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9608" agegroupid="7687" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7671" gender="M" number="34" order="13" round="FIN" preveventid="2082">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="9574" agegroupid="7672" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9575" agegroupid="7672" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7656" gender="F" number="31" order="8" round="FIN" preveventid="2034">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT heatid="9556" agegroupid="7657" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9557" agegroupid="7657" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7651" gender="M" number="30" order="9" round="FIN" preveventid="2027">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="9547" agegroupid="7652" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9548" agegroupid="7652" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2224" gender="F" number="41" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="2500" />
              <HEATS>
                <HEAT heatid="9618" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7681" gender="M" number="36" order="15" round="FIN" preveventid="5307">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="9600" agegroupid="7682" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9601" agegroupid="7682" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7641" gender="F" number="27" order="6" round="FIN" preveventid="2006">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT heatid="9532" agegroupid="7642" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9533" agegroupid="7642" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7666" gender="F" number="33" order="10" round="FIN" preveventid="2075">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT heatid="9568" agegroupid="7667" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9569" agegroupid="7667" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7631" gender="M" number="24" order="3" round="FIN" preveventid="1985">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="9517" agegroupid="7632" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9518" agegroupid="7632" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5333" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1062" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="5339" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="7676" gender="F" number="35" order="12" round="FIN" preveventid="2089">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="9589" agegroupid="7677" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9590" agegroupid="7677" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="2232" gender="M" number="42" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="2500" />
              <HEATS>
                <HEAT heatid="9619" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9620" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7626" gender="F" number="23" order="2" round="FIN" preveventid="1978">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="9507" agegroupid="7627" final="B" number="1" order="1" status="SEEDED" />
                <HEAT heatid="9508" agegroupid="7627" final="A" number="2" order="2" status="SEEDED" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1080" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1068" />
                <TIMESTANDARDREF marker="ENM" timestandardlistid="1072" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="4167" nation="GER" region="02" clubid="5520" name="1.SC Schweinfurt">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Severin" gender="M" lastname="Köhler" nation="GER" license="350064" athleteid="5521">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.55" entrycourse="SCM" eventid="1763" heatid="9378" lane="6">
                  <MEETINFO city="Lohr am Main" course="SCM" date="2019-03-24" name="Ufr.- &amp; 2. intern. Master-Kurzbahnmeisterschaften" qualificationtime="00:01:14.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.52" entrycourse="SCM" eventid="1985" heatid="9510" lane="4">
                  <MEETINFO city="Lohr am Main" course="SCM" date="2019-03-23" name="Ufr.- &amp; 2. intern. Master-Kurzbahnmeisterschaften" qualificationtime="00:00:33.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.37" entrycourse="SCM" eventid="1834" heatid="9446" lane="2">
                  <MEETINFO city="Lohr am Main" course="SCM" date="2019-03-24" name="Ufr.- &amp; 2. intern. Master-Kurzbahnmeisterschaften" qualificationtime="00:00:27.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.21" entrycourse="SCM" eventid="1971" heatid="9485" lane="5">
                  <MEETINFO city="Lohr am Main" course="SCM" date="2019-03-24" name="Ufr.- &amp; 2. intern. Master-Kurzbahnmeisterschaften" qualificationtime="00:00:59.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4224" nation="GER" region="02" clubid="5716" name="Delphin 77 Herzogenaurach">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Tim" gender="M" lastname="Dulitz" nation="GER" license="350454" athleteid="5717">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.25" entrycourse="SCM" eventid="1834" heatid="9450" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:25.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.12" entrycourse="SCM" eventid="1971" heatid="9494" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:55.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.63" entrycourse="LCM" eventid="5307" heatid="9592" lane="2">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:28.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Philipp" gender="M" lastname="Harig" nation="GER" license="300003" athleteid="5721">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.97" entrycourse="SCM" eventid="1749" heatid="9362" lane="5">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-12" name="Int. arena Swim Meeting" qualificationtime="00:02:04.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.63" entrycourse="SCM" eventid="1778" heatid="9393" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-05-25" name="18. Bamberg Open" qualificationtime="00:00:59.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.64" entrycourse="SCM" eventid="1971" heatid="9493" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-05-25" name="18. Bamberg Open" qualificationtime="00:00:55.64" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.92" entrycourse="SCM" eventid="2041" heatid="9559" lane="1">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:02:17.92" />
                </ENTRY>
                <ENTRY entrytime="00:04:24.93" entrycourse="SCM" eventid="2103" heatid="9611" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:24.93" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Xenia" gender="F" lastname="Schröder" nation="GER" license="415093" athleteid="5728">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.77" entrycourse="SCM" eventid="1756" heatid="9370" lane="6">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:36.77" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Sebastian" gender="M" lastname="Winkler" nation="GER" license="300000" athleteid="5730">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.44" entrycourse="SCM" eventid="1834" heatid="9453" lane="1">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:24.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.13" entrycourse="SCM" eventid="1971" heatid="9495" lane="5">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:54.09" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Paul" gender="M" lastname="Ziemainz" nation="GER" license="403946" athleteid="5733">
              <ENTRIES>
                <ENTRY entrytime="00:21:53.41" entrycourse="SCM" eventid="1792" heatid="9406" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:21:53.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4264" nation="GER" region="02" clubid="6901" name="MTV 1862 Pfaffenhofen/Ilm">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Hanna" gender="F" lastname="Schürer" nation="GER" license="328308" athleteid="6902">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.40" entrycourse="SCM" eventid="2089" heatid="9579" lane="4">
                  <MEETINFO city="Rain" course="SCM" date="2019-05-05" name="Tillystädter Schwimmen" qualificationtime="00:00:29.70" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="7077" nation="GER" region="02" clubid="5709" name="Nübad-Flipper">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Marie" gender="F" lastname="Brockhaus" nation="GER" license="199781" athleteid="5710">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.01" entrycourse="LCM" eventid="1059" heatid="9355" lane="3">
                  <MEETINFO city="Osnabrück" course="LCM" date="2019-02-24" name="15. schwimm-meeting Nettebad" qualificationtime="00:00:57.68" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.52" entrycourse="LCM" eventid="1785" heatid="9403" lane="3">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-05" name="69.Süddeutsche Meisterschaften" qualificationtime="00:01:05.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.21" entrycourse="LCM" eventid="1813" heatid="9426" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-04" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:02:13.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.01" entrycourse="LCM" eventid="1978" heatid="9506" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-03" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:02:03.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.83" entrycourse="LCM" eventid="2006" heatid="9531" lane="3">
                  <MEETINFO city="Heidelberg" course="LCM" date="2019-03-23" name="Nikar - Cup" qualificationtime="00:01:00.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4269" nation="GER" region="02" clubid="7691" name="Polizei SV Eichstätt">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Emanuel" gender="M" lastname="Höfl" nation="GER" license="256471" athleteid="7692">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.07" entrycourse="SCM" eventid="1834" heatid="9450" lane="3">
                  <MEETINFO city="Karlsruhe" course="LCM" date="2019-06-01" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:00:25.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.58" entrycourse="SCM" eventid="1971" heatid="9494" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:00:54.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.87" entrycourse="SCM" eventid="1985" heatid="9513" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:31.87" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Julia" gender="F" lastname="Iberle" nation="GER" license="313842" athleteid="7696">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.95" entrycourse="SCM" eventid="1059" heatid="9348" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:02.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.34" entrycourse="SCM" eventid="1799" heatid="9409" lane="2">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:13.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.89" entrycourse="SCM" eventid="2089" heatid="9582" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:28.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Florian" gender="M" lastname="Sattler" nation="GER" license="312155" athleteid="7700">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.71" entrycourse="SCM" eventid="1763" heatid="9381" lane="5">
                  <MEETINFO city="München" course="SCM" date="2019-05-12" name="24. Internationales Schwimmfest des MSV München" qualificationtime="00:01:09.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Magdalena" gender="F" lastname="Sattler" nation="GER" license="243094" athleteid="7702">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.46" entrycourse="SCM" eventid="1756" heatid="9373" lane="6">
                  <MEETINFO city="Karlsruhe" course="LCM" date="2019-06-01" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:00:35.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.83" entrycourse="SCM" eventid="1992" heatid="9522" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:17.83" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Jonas" gender="M" lastname="Schödl" nation="GER" license="329169" athleteid="7705">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.04" entrycourse="SCM" eventid="1763" heatid="9384" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:08.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.13" entrycourse="SCM" eventid="1985" heatid="9516" lane="1">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:31.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.92" entrycourse="SCM" eventid="2082" heatid="9572" lane="2">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:27.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="F" lastname="Vega Llamas" nation="GER" license="433387" athleteid="7709">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.89" entrycourse="SCM" eventid="1059" heatid="9346" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:05.40" />
                </ENTRY>
                <ENTRY entrytime="00:04:57.00" entrycourse="SCM" eventid="5320" heatid="9472" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:04:57.87" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.09" entrycourse="SCM" eventid="1978" heatid="9501" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:20.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.00" entrycourse="SCM" eventid="2089" heatid="9577" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:30.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4271" nation="GER" region="02" clubid="6604" name="Post-SV Nürnberg">
          <ATHLETES>
            <ATHLETE birthdate="2006-01-01" firstname="Artur" gender="M" lastname="Wölk" nation="GER" license="362630" athleteid="6605">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.04" entrycourse="SCM" eventid="1834" heatid="9443" lane="1">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:27.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4280" nation="GER" region="02" clubid="5553" name="SB Delphin 03 Augsburg">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Dreher" nation="GER" license="395983" athleteid="5554">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.41" entrycourse="SCM" eventid="1059" heatid="9350" lane="6">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:02.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.63" entrycourse="SCM" eventid="1841" heatid="9460" lane="5">
                  <MEETINFO city="Stadtbergen" course="SCM" date="2019-04-28" name="Stadtberger Mehrkampftag" qualificationtime="00:00:30.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.49" entrycourse="SCM" eventid="2089" heatid="9583" lane="3">
                  <MEETINFO city="Memmingen" course="SCM" date="2019-05-30" name="27. Internationales Memminger Mau Schwimmfest" qualificationtime="00:00:28.49" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Johanna" gender="F" lastname="Plail" nation="GER" license="316745" athleteid="5558">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.05" entrycourse="SCM" eventid="1799" heatid="9414" lane="6">
                  <MEETINFO city="Memmingen" course="SCM" date="2019-05-30" name="27. Internationales Memminger Mau Schwimmfest" qualificationtime="00:01:10.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.30" entrycourse="SCM" eventid="1827" heatid="9438" lane="4">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:45.30" />
                </ENTRY>
                <ENTRY entrytime="00:04:52.05" eventid="5320" heatid="9473" lane="1" />
                <ENTRY entrytime="00:02:12.83" entrycourse="SCM" eventid="1978" heatid="9505" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:12.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.96" entrycourse="SCM" eventid="1992" heatid="9523" lane="5">
                  <MEETINFO city="Memmingen" course="SCM" date="2019-05-30" name="27. Internationales Memminger Mau Schwimmfest" qualificationtime="00:01:16.96" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.40" entrycourse="SCM" eventid="2075" heatid="9567" lane="1">
                  <MEETINFO city="Stadtbergen" course="SCM" date="2019-04-28" name="Stadtberger Mehrkampftag" qualificationtime="00:02:30.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.18" entrycourse="SCM" eventid="2089" heatid="9580" lane="3">
                  <MEETINFO city="Memmingen" course="SCM" date="2019-05-30" name="27. Internationales Memminger Mau Schwimmfest" qualificationtime="00:00:29.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4290" nation="GER" region="02" clubid="6904" name="SC 53 Landshut">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Erlis" gender="M" lastname="Fazlija" nation="GER" license="331793" athleteid="6905">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.59" entrycourse="SCM" eventid="1749" heatid="9358" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:02:09.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.42" entrycourse="SCM" eventid="1806" heatid="9420" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:29.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.78" entrycourse="SCM" eventid="1848" heatid="9467" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:02:17.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.93" entrycourse="SCM" eventid="2013" heatid="9537" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:01:02.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.38" entrycourse="SCM" eventid="2027" heatid="9542" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:06.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Erza" gender="F" lastname="Fazlija" nation="GER" license="364830" athleteid="6911">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.75" entrycourse="SCM" eventid="1785" heatid="9398" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:12.75" />
                </ENTRY>
                <ENTRY entrytime="00:04:51.06" entrycourse="SCM" eventid="5320" heatid="9473" lane="5">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:04:51.06" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.10" entrycourse="SCM" eventid="1978" heatid="9502" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:17.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.82" entrycourse="SCM" eventid="2034" heatid="9550" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-30" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:00:33.82" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.41" entrycourse="SCM" eventid="2096" heatid="9604" lane="1">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:31.41" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Alexander" gender="M" lastname="Fuchs" nation="GER" license="284273" athleteid="6917">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.75" entrycourse="SCM" eventid="1749" heatid="9360" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:02:07.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.66" entrycourse="SCM" eventid="1971" heatid="9486" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:58.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Marieke" gender="F" lastname="Jacobs" nation="GER" license="335466" athleteid="6920">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.46" entrycourse="SCM" eventid="1756" heatid="9370" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-30" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:00:36.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.00" entrycourse="SCM" eventid="1827" heatid="9437" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-30" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:02:54.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.87" entrycourse="SCM" eventid="1992" heatid="9520" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:20.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.53" entrycourse="SCM" eventid="2089" heatid="9579" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:00:29.87" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Anna" gender="F" lastname="Karl" nation="GER" license="344913" athleteid="6925">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.36" entrycourse="SCM" eventid="1992" heatid="9520" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:20.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Hannah" gender="F" lastname="Köhnke" nation="GER" license="314299" athleteid="6927">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.64" entrycourse="SCM" eventid="1059" heatid="9347" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:03.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.18" entrycourse="SCM" eventid="1785" heatid="9401" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:01:08.78" />
                </ENTRY>
                <ENTRY entrytime="00:04:49.70" entrycourse="LCM" eventid="5320" heatid="9473" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:49.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.29" entrycourse="SCM" eventid="1978" heatid="9503" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:02:16.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.72" entrycourse="SCM" eventid="2006" heatid="9529" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-30" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:01:08.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.89" entrycourse="SCM" eventid="2034" heatid="9552" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-30" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:00:32.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.55" entrycourse="SCM" eventid="2096" heatid="9604" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:02:27.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Daniel" gender="M" lastname="Siminenko" nation="GER" license="300185" athleteid="6935">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.20" entrycourse="SCM" eventid="1763" heatid="9384" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:07.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.99" entrycourse="SCM" eventid="1778" heatid="9391" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:00.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.96" entrycourse="SCM" eventid="1834" heatid="9451" lane="5">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:25.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.44" entrycourse="SCM" eventid="1985" heatid="9516" lane="6">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:31.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.85" entrycourse="SCM" eventid="2027" heatid="9545" lane="2">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:01.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.17" entrycourse="SCM" eventid="5307" heatid="9595" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:27.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4286" nation="GER" region="02" clubid="5566" name="SC Delphin Ingolstadt">
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Jonas" gender="M" lastname="Drieling" nation="GER" license="280053" athleteid="5567">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.40" entrycourse="SCM" eventid="1806" heatid="9422" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:26.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.40" eventid="1834" heatid="9452" lane="5" />
                <ENTRY entrytime="00:01:00.50" eventid="2013" heatid="9538" lane="2" />
                <ENTRY entrytime="00:00:25.80" eventid="5307" heatid="9599" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Maximilian" gender="M" lastname="Hagl" nation="GER" license="341127" athleteid="5572">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.75" entrycourse="SCM" eventid="1749" heatid="9360" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:05.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.40" entrycourse="SCM" eventid="1806" heatid="9422" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:29.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.00" entrycourse="SCM" eventid="1848" heatid="9468" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:20.12" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.80" entrycourse="SCM" eventid="2013" heatid="9535" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:03.76" />
                </ENTRY>
                <ENTRY entrytime="00:04:28.00" entrycourse="SCM" eventid="2103" heatid="9611" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:28.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Fabian" gender="M" lastname="Heinemann" nation="GER" license="313851" athleteid="5578">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.80" entrycourse="SCM" eventid="1778" heatid="9394" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:59.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.10" entrycourse="SCM" eventid="1806" heatid="9420" lane="2">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:27.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.20" entrycourse="SCM" eventid="1834" heatid="9454" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:24.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.90" entrycourse="SCM" eventid="1971" heatid="9497" lane="5">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:52.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.60" entrycourse="SCM" eventid="2027" heatid="9545" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:00.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.20" entrycourse="SCM" eventid="5307" heatid="9599" lane="5">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:26.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Larissa" gender="F" lastname="Heinemann" nation="GER" license="313844" athleteid="5585">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" entrycourse="SCM" eventid="1059" heatid="9354" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:00.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.20" entrycourse="SCM" eventid="1799" heatid="9414" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:07.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.80" entrycourse="SCM" eventid="1841" heatid="9461" lane="2">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-03" name="69.Süddeutsche Meisterschaften" qualificationtime="00:00:29.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.60" entrycourse="SCM" eventid="2006" heatid="9530" lane="2">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-05" name="69.Süddeutsche Meisterschaften" qualificationtime="00:01:06.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.90" entrycourse="SCM" eventid="2089" heatid="9586" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:27.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Joshua" gender="M" lastname="Hollweck" nation="GER" license="313850" athleteid="5593">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.40" entrycourse="SCM" eventid="1778" heatid="9394" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:00.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.40" entrycourse="SCM" eventid="1820" heatid="9431" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:16.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.60" entrycourse="LCM" eventid="1834" heatid="9449" lane="1">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-05" name="69.Süddeutsche Meisterschaften" qualificationtime="00:00:26.05" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.40" entrycourse="SCM" eventid="1971" heatid="9493" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:56.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.20" eventid="2027" heatid="9545" lane="5" />
                <ENTRY entrytime="00:00:27.20" entrycourse="LCM" eventid="5307" heatid="9595" lane="2">
                  <MEETINFO city="Pfaffenhofen" course="LCM" date="2019-06-30" name="Kreispokal  Kreis V Obb." qualificationtime="00:00:27.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Valerie" gender="F" lastname="Höfl" nation="GER" license="363083" athleteid="5591">
              <ENTRIES>
                <ENTRY entrytime="00:02:55.40" entrycourse="SCM" eventid="1827" heatid="9436" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:54.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Maria" gender="F" lastname="Kapfer" nation="GER" license="322566" athleteid="5600">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.50" entrycourse="SCM" eventid="1785" heatid="9403" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:07.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.20" entrycourse="SCM" eventid="1799" heatid="9415" lane="5">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-10" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:01:09.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.50" entrycourse="SCM" eventid="1827" heatid="9439" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:02:45.37" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.00" entrycourse="SCM" eventid="1978" heatid="9506" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:13.56" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.00" entrycourse="SCM" eventid="2075" heatid="9566" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:02:29.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.80" entrycourse="SCM" eventid="2096" heatid="9605" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:25.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Ariana" gender="F" lastname="Lind" nation="GER" license="356602" athleteid="5607">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.88" entrycourse="SCM" eventid="2089" heatid="9578" lane="2">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:29.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Claudius" gender="M" lastname="Lindner" nation="GER" license="331306" athleteid="5609">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.65" entrycourse="SCM" eventid="1806" heatid="9422" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:28.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.60" entrycourse="SCM" eventid="1834" heatid="9445" lane="6">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:26.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.50" entrycourse="SCM" eventid="1848" heatid="9468" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:17.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.40" entrycourse="SCM" eventid="1971" heatid="9487" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:58.90" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.00" entrycourse="SCM" eventid="2013" heatid="9536" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:03.05" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.80" entrycourse="SCM" eventid="5307" heatid="9591" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:28.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Katharina" gender="F" lastname="Marb" nation="GER" license="300191" athleteid="5616">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.50" entrycourse="SCM" eventid="1059" heatid="9355" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:00.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.50" entrycourse="SCM" eventid="1785" heatid="9403" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:05.51" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.80" entrycourse="SCM" eventid="1978" heatid="9506" lane="5">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-09" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:02:12.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.40" entrycourse="SCM" eventid="2034" heatid="9554" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:30.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.80" entrycourse="SCM" eventid="2096" heatid="9605" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:22.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Leonie" gender="F" lastname="Mathe" nation="GER" license="215384" athleteid="5622">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.30" entrycourse="SCM" eventid="1059" heatid="9355" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:00:57.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.60" entrycourse="SCM" eventid="1756" heatid="9373" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:33.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.00" entrycourse="SCM" eventid="1992" heatid="9524" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:12.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.00" entrycourse="SCM" eventid="2089" heatid="9588" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:00:26.72" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Christoph" gender="M" lastname="Mooser" nation="GER" license="240870" athleteid="5627">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" entrycourse="SCM" eventid="1763" heatid="9383" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:05.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.60" entrycourse="SCM" eventid="1806" heatid="9421" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:27.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.80" entrycourse="SCM" eventid="1985" heatid="9514" lane="3">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-10" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:00:29.34" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.20" entrycourse="SCM" eventid="2027" heatid="9544" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:59.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.00" entrycourse="SCM" eventid="2082" heatid="9572" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:20.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Debora" gender="F" lastname="Mooser" nation="GER" license="334714" athleteid="5633">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.94" entrycourse="SCM" eventid="1756" heatid="9369" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:36.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.08" entrycourse="SCM" eventid="1992" heatid="9519" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:21.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.95" entrycourse="SCM" eventid="2089" heatid="9577" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:29.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Emely" gender="F" lastname="Neumüller" nation="GER" license="352380" athleteid="5637">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.00" entrycourse="SCM" eventid="1059" heatid="9348" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:03.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.80" entrycourse="SCM" eventid="1785" heatid="9398" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:12.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.65" entrycourse="SCM" eventid="1841" heatid="9460" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:30.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.60" entrycourse="SCM" eventid="2034" heatid="9551" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:33.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.95" entrycourse="SCM" eventid="2089" heatid="9582" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:28.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Isabell" gender="F" lastname="Schiller" nation="GER" license="322565" athleteid="5643">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.20" entrycourse="SCM" eventid="1785" heatid="9403" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:07.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.60" eventid="1799" heatid="9412" lane="2" />
                <ENTRY entrytime="00:00:30.80" entrycourse="SCM" eventid="1841" heatid="9459" lane="2">
                  <MEETINFO city="Pfaffenhofen" course="LCM" date="2019-06-30" name="Kreispokal  Kreis V Obb." qualificationtime="00:00:30.06" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.20" entrycourse="SCM" eventid="1992" heatid="9524" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:17.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.90" entrycourse="SCM" eventid="2075" heatid="9565" lane="2">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-09" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:02:27.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.80" entrycourse="SCM" eventid="2096" heatid="9606" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:23.24" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Johanna" gender="F" lastname="Schmid" nation="GER" license="266871" athleteid="5650">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.12" entrycourse="SCM" eventid="1756" heatid="9373" lane="5">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:36.19" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Christina" gender="F" lastname="Schulz" nation="GER" license="352365" athleteid="5652">
              <ENTRIES>
                <ENTRY entrytime="00:02:51.80" entrycourse="SCM" eventid="1827" heatid="9439" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:50.25" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.80" entrycourse="SCM" eventid="1978" heatid="9500" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:20.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Josy Cindy" gender="F" lastname="Urban" nation="GER" license="345861" athleteid="5655">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.83" entrycourse="SCM" eventid="1756" heatid="9369" lane="3">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-10" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:00:36.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.14" entrycourse="SCM" eventid="2089" heatid="9581" lane="2">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-05" name="69.Süddeutsche Meisterschaften" qualificationtime="00:00:29.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Emma Johanna" gender="F" lastname="Weiß" nation="GER" license="317378" athleteid="5658">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.80" entrycourse="SCM" eventid="1756" heatid="9372" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:33.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.00" eventid="1799" heatid="9413" lane="2" />
                <ENTRY entrytime="00:00:31.20" entrycourse="SCM" eventid="1841" heatid="9458" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:31.18" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.60" entrycourse="SCM" eventid="1992" heatid="9524" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:16.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.80" entrycourse="SCM" eventid="2034" heatid="9554" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:31.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.20" entrycourse="SCM" eventid="2089" heatid="9587" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:00:27.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.40" eventid="5316" heatid="9481" lane="4" />
                <ENTRY entrytime="00:01:38.40" eventid="2232" heatid="9620" lane="2" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.00" eventid="5314" heatid="9483" lane="5">
                  <MEETINFO city="Karlsruhe" date="2019-05-31" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:02:23.89" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.80" eventid="2224" heatid="9618" lane="2">
                  <MEETINFO city="Karlsruhe" date="2019-05-31" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:02:08.02" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:42.60" eventid="1855" heatid="9477" lane="4">
                  <MEETINFO city="Erding" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:34.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.40" eventid="5303" heatid="9615" lane="2">
                  <MEETINFO city="Pfaffenhofen" date="2019-06-30" name="Kreispokal  Kreis V Obb." qualificationtime="00:02:01.20" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4292" nation="GER" region="02" clubid="6607" name="SC Prinz Eugen München">
          <ATHLETES>
            <ATHLETE birthdate="2006-01-01" firstname="Johanna" gender="F" lastname="Berger" nation="GER" license="361332" athleteid="6608">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.86" entrycourse="SCM" eventid="1059" heatid="9349" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:01:02.86" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.91" entrycourse="SCM" eventid="1756" heatid="9371" lane="2">
                  <MEETINFO city="Neufahrn" course="SCM" date="2019-07-13" name="Neufahrner Pokalschwimmen" qualificationtime="00:00:35.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.07" entrycourse="SCM" eventid="1799" heatid="9410" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:12.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.46" entrycourse="SCM" eventid="1841" heatid="9458" lane="6">
                  <MEETINFO city="Wetzlar" course="LCM" date="2019-05-05" name="27. Süddeutsche Jahrgangsmeisterschaften" qualificationtime="00:00:31.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.12" entrycourse="SCM" eventid="1992" heatid="9521" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:01:19.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.74" entrycourse="SCM" eventid="2089" heatid="9583" lane="1">
                  <MEETINFO city="Wetzlar" course="LCM" date="2019-05-04" name="27. Süddeutsche Jahrgangsmeisterschaften" qualificationtime="00:00:28.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Hanna" gender="F" lastname="Pfannes" nation="GER" license="301469" athleteid="6615">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.57" entrycourse="SCM" eventid="1756" heatid="9372" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:34.66" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.53" entrycourse="SCM" eventid="1785" heatid="9402" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:06.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.62" entrycourse="SCM" eventid="1827" heatid="9438" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:37.62" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.09" entrycourse="SCM" eventid="1992" heatid="9522" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:15.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.52" entrycourse="SCM" eventid="2034" heatid="9555" lane="4">
                  <MEETINFO city="Neufahrn" course="SCM" date="2019-07-13" name="Neufahrner Pokalschwimmen" qualificationtime="00:00:30.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Maya" gender="F" lastname="Rainer" nation="GER" license="339440" athleteid="6621">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.98" entrycourse="SCM" eventid="1059" heatid="9353" lane="2">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-17" name="10. Internationales Frühjahresmeeting" qualificationtime="00:00:59.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.92" entrycourse="SCM" eventid="1785" heatid="9401" lane="4">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-16" name="10. Internationales Frühjahresmeeting" qualificationtime="00:01:06.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.63" entrycourse="SCM" eventid="1799" heatid="9412" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:10.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.26" entrycourse="SCM" eventid="2089" heatid="9586" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:26.27" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Maria" gender="F" lastname="Vollmer" nation="GER" license="297327" athleteid="6626">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.11" entrycourse="SCM" eventid="1059" heatid="9352" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:01:01.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.77" entrycourse="SCM" eventid="1756" heatid="9371" lane="4">
                  <MEETINFO city="München Obergiesing" course="SCM" date="2019-03-23" name="OMP Frühjahrsdurchgang - Offen/Minis" qualificationtime="00:00:36.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:46.83" entrycourse="SCM" eventid="1827" heatid="9438" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:46.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.59" entrycourse="SCM" eventid="1978" heatid="9503" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:15.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.52" entrycourse="SCM" eventid="1992" heatid="9524" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:01:17.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.78" entrycourse="SCM" eventid="2075" heatid="9564" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:32.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.14" entrycourse="SCM" eventid="2089" heatid="9585" lane="6">
                  <MEETINFO city="München Obergiesing" course="SCM" date="2019-03-23" name="OMP Frühjahrsdurchgang - Offen/Minis" qualificationtime="00:00:28.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.43" eventid="5314" heatid="9483" lane="2">
                  <MEETINFO city="München Obergiesing" date="2019-03-23" name="OMP Frühjahrsdurchgang - Offen/Minis" qualificationtime="00:02:13.08" />
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6615" number="1" />
                    <RELAYPOSITION athleteid="6608" number="2" />
                    <RELAYPOSITION athleteid="6626" number="3" />
                    <RELAYPOSITION athleteid="6621" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:53.34" eventid="2224" heatid="9618" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6621" number="1" />
                    <RELAYPOSITION athleteid="6608" number="2" />
                    <RELAYPOSITION athleteid="6615" number="3" />
                    <RELAYPOSITION athleteid="6626" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6524" nation="GER" region="02" clubid="6493" name="SC Regensburg">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Ines" gender="F" lastname="Erban" nation="GER" license="343982" athleteid="6494">
              <ENTRIES>
                <ENTRY entrytime="00:04:49.00" entrycourse="SCM" eventid="5320" heatid="9473" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:43.34" />
                </ENTRY>
                <ENTRY entrytime="00:18:38.91" entrycourse="LCM" eventid="5318" heatid="9479" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:18:38.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Jakob" gender="M" lastname="Erban" nation="GER" license="333295" athleteid="6497">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.26" entrycourse="SCM" eventid="1749" heatid="9362" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:02:03.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.70" entrycourse="LCM" eventid="1834" heatid="9444" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:26.96" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lena" gender="F" lastname="Gerl" nation="GER" license="370044" athleteid="6500">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.04" entrycourse="SCM" eventid="1059" heatid="9345" lane="3">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:04.92" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.03" entrycourse="SCM" eventid="1813" heatid="9425" lane="1">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:36.03" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.27" entrycourse="SCM" eventid="1978" heatid="9501" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:19.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.62" entrycourse="SCM" eventid="2075" heatid="9562" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:36.11" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Leon" gender="M" lastname="Heberlein" nation="GER" license="336955" athleteid="6505">
              <ENTRIES>
                <ENTRY entrytime="00:02:08.63" entrycourse="SCM" eventid="1749" heatid="9359" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:08.63" />
                </ENTRY>
                <ENTRY entrytime="00:17:44.03" entrycourse="SCM" eventid="1792" heatid="9407" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:17:44.03" />
                </ENTRY>
                <ENTRY entrytime="00:04:29.26" entrycourse="LCM" eventid="2103" heatid="9610" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:29.26" />
                </ENTRY>
                <ENTRY entrytime="00:09:16.48" entrycourse="LCM" eventid="2168" heatid="9616" lane="5">
                  <MEETINFO city="Graz-Eggenberg" course="LCM" date="2019-04-28" name="Int. Ströck ATUS Graz Trophy" qualificationtime="00:09:16.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Alexandra" gender="F" lastname="Jaud" nation="GER" license="332959" athleteid="6510">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.28" entrycourse="SCM" eventid="1756" heatid="9369" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:37.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.32" entrycourse="SCM" eventid="1799" heatid="9409" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:13.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.22" entrycourse="LCM" eventid="1827" heatid="9436" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:56.22" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.60" entrycourse="SCM" eventid="1992" heatid="9520" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:19.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.12" entrycourse="SCM" eventid="2075" heatid="9563" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:36.07" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Anne" gender="F" lastname="Mauerer" nation="GER" license="299448" athleteid="6516">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.00" entrycourse="SCM" eventid="1059" heatid="9350" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:01:01.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.16" entrycourse="SCM" eventid="1756" heatid="9374" lane="1">
                  <MEETINFO city="Magdeburg" course="LCM" date="2019-03-30" name="29. Pokal der Gothaer Versicherung" qualificationtime="00:00:35.16" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.42" entrycourse="SCM" eventid="1785" heatid="9401" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:07.37" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.50" entrycourse="SCM" eventid="1799" heatid="9415" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:07.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:49.50" entrycourse="LCM" eventid="1827" heatid="9437" lane="5">
                  <MEETINFO city="Magdeburg" course="LCM" date="2019-03-30" name="29. Pokal der Gothaer Versicherung" qualificationtime="00:02:45.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.20" entrycourse="SCM" eventid="1841" heatid="9461" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:29.75" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.29" entrycourse="SCM" eventid="1978" heatid="9504" lane="6">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-07" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:02:11.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.50" entrycourse="SCM" eventid="1992" heatid="9522" lane="1">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-17" name="10. Internationales Frühjahresmeeting" qualificationtime="00:01:16.58" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.00" entrycourse="SCM" eventid="2006" heatid="9528" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:07.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.90" entrycourse="SCM" eventid="2034" heatid="9555" lane="5">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:31.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.00" entrycourse="SCM" eventid="2075" heatid="9565" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-07" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:02:27.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Justus" gender="M" lastname="Menzel" nation="GER" license="336910" athleteid="6528">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.60" entrycourse="SCM" eventid="1749" heatid="9358" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:09.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.60" entrycourse="SCM" eventid="1806" heatid="9419" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:29.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.05" entrycourse="SCM" eventid="1834" heatid="9443" lane="6">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:26.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.71" entrycourse="SCM" eventid="1848" heatid="9467" lane="1">
                  <MEETINFO city="Parsberg" course="SCM" date="2019-02-24" name="DMS  Bezirksliga" qualificationtime="00:02:18.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.96" entrycourse="SCM" eventid="1971" heatid="9485" lane="4">
                  <MEETINFO city="Parsberg" course="SCM" date="2019-02-24" name="DMS  Bezirksliga" qualificationtime="00:00:59.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.75" entrycourse="SCM" eventid="2013" heatid="9535" lane="5">
                  <MEETINFO city="Parsberg" course="SCM" date="2019-02-24" name="DMS  Bezirksliga" qualificationtime="00:01:04.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Alexander" gender="M" lastname="Metzler" nation="GER" license="305951" athleteid="6535">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.26" entrycourse="SCM" eventid="1749" heatid="9365" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:54.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.83" entrycourse="SCM" eventid="1763" heatid="9381" lane="1">
                  <MEETINFO city="Magdeburg" course="LCM" date="2019-03-31" name="29. Pokal der Gothaer Versicherung" qualificationtime="00:01:09.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.23" entrycourse="SCM" eventid="1778" heatid="9392" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:59.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.76" entrycourse="SCM" eventid="1806" heatid="9421" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:27.57" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.43" entrycourse="SCM" eventid="1820" heatid="9433" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:11.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.60" entrycourse="SCM" eventid="1834" heatid="9449" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:25.26" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.90" entrycourse="SCM" eventid="1848" heatid="9469" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:11.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.17" entrycourse="SCM" eventid="1971" heatid="9492" lane="5">
                  <MEETINFO city="Magdeburg" course="LCM" date="2019-03-30" name="29. Pokal der Gothaer Versicherung" qualificationtime="00:00:56.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.49" entrycourse="SCM" eventid="1985" heatid="9512" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:31.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.59" entrycourse="SCM" eventid="2013" heatid="9537" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:59.45" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.55" entrycourse="SCM" eventid="2027" heatid="9546" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:01.02" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.26" entrycourse="LCM" eventid="2082" heatid="9573" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-16" name="10. Internationales Frühjahresmeeting" qualificationtime="00:02:30.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.07" entrycourse="SCM" eventid="5307" heatid="9596" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:27.04" />
                </ENTRY>
                <ENTRY entrytime="00:04:15.61" entrycourse="LCM" eventid="2103" heatid="9612" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:04:15.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Michael" gender="M" lastname="Moser" nation="GER" license="356878" athleteid="6550">
              <ENTRIES>
                <ENTRY entrytime="00:02:08.36" entrycourse="SCM" eventid="1749" heatid="9359" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:08.36" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.40" entrycourse="SCM" eventid="1778" heatid="9390" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:01:02.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.70" entrycourse="SCM" eventid="1820" heatid="9430" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:24.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.83" entrycourse="SCM" eventid="2041" heatid="9559" lane="6">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:02:22.83" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Mark" gender="M" lastname="Nickles" nation="GER" license="309205" athleteid="6555">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.08" entrycourse="SCM" eventid="1778" heatid="9391" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:01.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.60" entrycourse="SCM" eventid="1806" heatid="9421" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:28.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.01" entrycourse="SCM" eventid="1834" heatid="9448" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:26.01" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.19" entrycourse="SCM" eventid="1848" heatid="9469" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:17.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.50" entrycourse="SCM" eventid="1985" heatid="9512" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:32.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.39" entrycourse="SCM" eventid="2013" heatid="9538" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:01:02.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.70" entrycourse="SCM" eventid="5307" heatid="9594" lane="4">
                  <MEETINFO city="Graz-Eggenberg" course="LCM" date="2019-04-28" name="Int. Ströck ATUS Graz Trophy" qualificationtime="00:00:27.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Tiffany Vanessa" gender="F" lastname="Salva" nation="GER" license="331446" athleteid="6563">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.02" entrycourse="SCM" eventid="1059" heatid="9348" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:03.02" />
                </ENTRY>
                <ENTRY entrytime="00:05:32.04" entrycourse="LCM" eventid="1771" heatid="9387" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-01-19" name="Bayerische Meisterschaften lange Strecken" qualificationtime="00:05:32.04" />
                </ENTRY>
                <ENTRY entrytime="00:04:43.23" entrycourse="SCM" eventid="5320" heatid="9474" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:04:43.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.67" entrycourse="LCM" eventid="1978" heatid="9502" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:17.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Elisabeth" gender="F" lastname="Striepling" nation="GER" license="307177" athleteid="6568">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.35" entrycourse="SCM" eventid="1799" heatid="9412" lane="3">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:12.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.42" entrycourse="SCM" eventid="1841" heatid="9460" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:29.18" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.87" entrycourse="SCM" eventid="2006" heatid="9531" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:06.87" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.10" entrycourse="SCM" eventid="2075" heatid="9564" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:31.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.50" entrycourse="SCM" eventid="2089" heatid="9583" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:28.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Robin" gender="M" lastname="Swoboda" nation="GER" license="279876" athleteid="6574">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.17" entrycourse="SCM" eventid="1749" heatid="9360" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:05.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.02" entrycourse="SCM" eventid="1763" heatid="9379" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:11.01" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.00" entrycourse="SCM" eventid="1778" heatid="9389" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:02.95" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.43" entrycourse="SCM" eventid="1834" heatid="9446" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:26.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.02" entrycourse="SCM" eventid="1971" heatid="9488" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:57.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.33" entrycourse="SCM" eventid="1985" heatid="9512" lane="3">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:31.77" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.59" entrycourse="SCM" eventid="2027" heatid="9543" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:01:04.59" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.82" entrycourse="SCM" eventid="2082" heatid="9571" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:35.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.49" entrycourse="SCM" eventid="5307" heatid="9592" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:28.49" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Amira" gender="F" lastname="Varna" nation="GER" license="358238" athleteid="6584">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.55" entrycourse="SCM" eventid="1059" heatid="9347" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:03.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.77" entrycourse="SCM" eventid="1785" heatid="9398" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:12.77" />
                </ENTRY>
                <ENTRY entrytime="00:04:54.00" entrycourse="LCM" eventid="5320" heatid="9473" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:52.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.12" entrycourse="SCM" eventid="1978" heatid="9501" lane="3">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-12" name="Int. arena Swim Meeting" qualificationtime="00:02:19.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.90" entrycourse="SCM" eventid="2034" heatid="9550" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:33.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.27" entrycourse="SCM" eventid="2089" heatid="9576" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:29.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.00" entrycourse="SCM" eventid="2096" heatid="9602" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:35.76" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Nele" gender="F" lastname="Weinfurtner" nation="GER" license="260402" athleteid="6592">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.68" entrycourse="SCM" eventid="1756" heatid="9372" lane="6">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:00:35.53" />
                </ENTRY>
                <ENTRY entrytime="00:05:10.39" entrycourse="LCM" eventid="1771" heatid="9388" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:05:12.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.30" entrycourse="SCM" eventid="1785" heatid="9402" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:07.39" />
                </ENTRY>
                <ENTRY entrytime="00:04:38.00" entrycourse="SCM" eventid="5320" heatid="9475" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:37.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.10" entrycourse="SCM" eventid="1978" heatid="9506" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:11.10" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.95" entrycourse="SCM" eventid="2075" heatid="9565" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:02:25.95" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.50" entrycourse="SCM" eventid="2096" heatid="9604" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:20.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.07" eventid="5316" heatid="9481" lane="6">
                  <MEETINFO city="Dachau" date="2019-02-16" name="20. Int. Dachauer Masters-Cup" qualificationtime="00:02:03.27" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.31" eventid="5314" heatid="9482" lane="3">
                  <MEETINFO city="Dachau" date="2019-02-16" name="20. Int. Dachauer Masters-Cup" qualificationtime="00:02:30.42" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.00" eventid="1855" heatid="9476" lane="3">
                  <MEETINFO city="Dachau" date="2019-02-17" name="20. Int. Dachauer Masters-Cup" qualificationtime="00:02:10.67" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.00" eventid="5303" heatid="9614" lane="4">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:02:09.26" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4296" nation="GER" region="02" clubid="6958" name="SC Wfr. München">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Johanna" gender="F" lastname="Bander" nation="GER" license="281505" athleteid="6959">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.46" entrycourse="SCM" eventid="1059" heatid="9349" lane="4">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:01:02.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.41" entrycourse="LCM" eventid="1841" heatid="9458" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:30.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.46" entrycourse="SCM" eventid="2006" heatid="9528" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:09.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.66" entrycourse="SCM" eventid="2089" heatid="9583" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:28.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Alexander" gender="M" lastname="Bender" nation="GER" license="323184" athleteid="6964">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.25" entrycourse="SCM" eventid="1763" heatid="9379" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:11.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.23" entrycourse="SCM" eventid="1985" heatid="9510" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:33.24" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Stella" gender="F" lastname="Da Silva Buttkus" nation="GER" license="384713" athleteid="6967">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.87" entrycourse="SCM" eventid="1059" heatid="9347" lane="6">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:03.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.25" entrycourse="SCM" eventid="2089" heatid="9580" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:29.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Paul" gender="M" lastname="Deuker" nation="GER" license="248532" athleteid="6970">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.82" entrycourse="SCM" eventid="1778" heatid="9393" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:58.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.72" entrycourse="SCM" eventid="1834" heatid="9453" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:24.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.79" entrycourse="SCM" eventid="1971" heatid="9496" lane="1">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-09" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:00:54.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.44" entrycourse="SCM" eventid="5307" heatid="9598" lane="5">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-09" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:00:27.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Alexander" gender="M" lastname="Gubanov" nation="GER" license="243921" athleteid="6978">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.32" entrycourse="SCM" eventid="1763" heatid="9381" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:09.69" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Michael" gender="M" lastname="Gubanov" nation="GER" license="261412" athleteid="6980">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.44" entrycourse="SCM" eventid="1834" heatid="9449" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:00:25.44" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Greta" gender="F" lastname="Heinzelmann" nation="GER" license="173466" athleteid="6982">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.54" entrycourse="SCM" eventid="1059" heatid="9353" lane="4">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-01-12" name="34. Augsburger Zirbelnuss-Schwimmen" qualificationtime="00:01:02.16" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.68" entrycourse="SCM" eventid="1785" heatid="9402" lane="4">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-01-13" name="34. Augsburger Zirbelnuss-Schwimmen" qualificationtime="00:01:09.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.95" entrycourse="SCM" eventid="2034" heatid="9555" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:30.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.96" entrycourse="SCM" eventid="2089" heatid="9587" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:27.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Oliver" gender="M" lastname="Hoffmann" nation="GER" license="270010" athleteid="6987">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.99" entrycourse="SCM" eventid="1763" heatid="9384" lane="2">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-01-12" name="34. Augsburger Zirbelnuss-Schwimmen" qualificationtime="00:01:07.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.66" entrycourse="SCM" eventid="1806" heatid="9420" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:27.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.08" entrycourse="SCM" eventid="1848" heatid="9467" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:09.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.81" entrycourse="SCM" eventid="1985" heatid="9515" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:30.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.67" entrycourse="SCM" eventid="2013" heatid="9536" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-01-13" name="34. Augsburger Zirbelnuss-Schwimmen" qualificationtime="00:00:58.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.80" entrycourse="SCM" eventid="5307" heatid="9598" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:26.80" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Jamie" gender="M" lastname="Holmes" nation="GER" license="330605" athleteid="6994">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.60" entrycourse="SCM" eventid="1749" heatid="9358" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:09.46" />
                </ENTRY>
                <ENTRY entrytime="00:18:07.23" entrycourse="LCM" eventid="1792" heatid="9406" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-02-23" name="30. Süddeutsche Meisterschaften Lange Strecken" qualificationtime="00:18:07.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.92" entrycourse="SCM" eventid="1971" heatid="9485" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:58.07" />
                </ENTRY>
                <ENTRY entrytime="00:04:32.63" entrycourse="SCM" eventid="2103" heatid="9610" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:04:26.96" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Nate" gender="M" lastname="Holmes" nation="GER" license="335037" athleteid="6999">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.42" entrycourse="SCM" eventid="1749" heatid="9359" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:09.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.86" entrycourse="SCM" eventid="1763" heatid="9377" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:14.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.02" entrycourse="SCM" eventid="1820" heatid="9430" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:25.02" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.35" entrycourse="SCM" eventid="1848" heatid="9466" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:24.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.81" entrycourse="SCM" eventid="1971" heatid="9486" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:58.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.19" entrycourse="SCM" eventid="1985" heatid="9509" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:34.19" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.53" entrycourse="SCM" eventid="2013" heatid="9534" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:06.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Moritz" gender="M" lastname="Kolmberger" nation="GER" license="369011" athleteid="7010">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.04" entrycourse="SCM" eventid="1749" heatid="9362" lane="1">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:04.04" />
                </ENTRY>
                <ENTRY entrytime="00:17:57.47" entrycourse="SCM" eventid="1792" heatid="9406" lane="3">
                  <MEETINFO city="Rosenheim" course="LCM" date="2019-05-31" name="30. Int. Langstreckenschwimmen" qualificationtime="00:17:57.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.18" entrycourse="SCM" eventid="1834" heatid="9442" lane="4">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:00:26.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.02" entrycourse="SCM" eventid="1971" heatid="9488" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:58.01" />
                </ENTRY>
                <ENTRY entrytime="00:04:25.82" entrycourse="SCM" eventid="2103" heatid="9611" lane="2">
                  <MEETINFO city="Rosenheim" course="LCM" date="2019-06-02" name="30. Int. Langstreckenschwimmen" qualificationtime="00:04:25.82" />
                </ENTRY>
                <ENTRY entrytime="00:09:15.34" entrycourse="LCM" eventid="2168" heatid="9616" lane="2">
                  <MEETINFO city="Rosenheim" course="LCM" date="2019-06-01" name="30. Int. Langstreckenschwimmen" qualificationtime="00:09:15.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Nicolas" gender="M" lastname="Kolmberger" nation="GER" license="369012" athleteid="7017">
              <ENTRIES>
                <ENTRY entrytime="00:18:36.37" entrycourse="SCM" eventid="1792" heatid="9406" lane="5">
                  <MEETINFO city="Bad Tölz" course="SCM" date="2019-02-24" name="DMS Bezirksdurchgang Oberbayern" qualificationtime="00:18:36.37" />
                </ENTRY>
                <ENTRY entrytime="00:09:55.03" entrycourse="LCM" eventid="2168" status="RJC">
                  <MEETINFO city="Rosenheim" course="LCM" date="2019-06-01" name="30. Int. Langstreckenschwimmen" qualificationtime="00:09:55.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Paul" gender="M" lastname="Melcer" nation="GER" license="296353" athleteid="7020">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.55" entrycourse="SCM" eventid="1806" heatid="9422" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:28.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.50" entrycourse="SCM" eventid="1834" heatid="9445" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:26.38" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.00" entrycourse="SCM" eventid="1848" heatid="9467" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:14.67" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.75" entrycourse="SCM" eventid="1971" heatid="9486" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:57.71" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.42" entrycourse="SCM" eventid="2013" heatid="9537" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:01.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.06" entrycourse="SCM" eventid="2027" heatid="9545" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:04.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Daniil" gender="M" lastname="Melnik" nation="GER" license="269642" athleteid="7027">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.80" entrycourse="SCM" eventid="1985" heatid="9514" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:31.85" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Rachel" gender="F" lastname="Omoruyi" nation="GER" license="302750" athleteid="7032">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.42" entrycourse="SCM" eventid="1059" heatid="9349" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:02.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.80" entrycourse="SCM" eventid="1785" heatid="9399" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:11.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.39" entrycourse="SCM" eventid="1799" heatid="9411" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:10.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.13" entrycourse="SCM" eventid="1978" heatid="9502" lane="4">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-12" name="Int. arena Swim Meeting" qualificationtime="00:02:17.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.26" entrycourse="SCM" eventid="2089" heatid="9584" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:28.26" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.30" entrycourse="LCM" eventid="2096" heatid="9604" lane="6">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-12" name="Int. arena Swim Meeting" qualificationtime="00:02:34.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Esther" gender="F" lastname="Pearce" nation="GER" license="394966" athleteid="7039">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.03" entrycourse="SCM" eventid="1756" heatid="9371" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-16" name="10. Internationales Frühjahresmeeting" qualificationtime="00:00:36.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.48" entrycourse="SCM" eventid="1799" heatid="9410" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:12.48" />
                </ENTRY>
                <ENTRY entrytime="00:02:46.28" entrycourse="SCM" eventid="1827" heatid="9439" lane="2">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:46.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.00" entrycourse="SCM" eventid="1992" heatid="9521" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:18.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.16" entrycourse="SCM" eventid="2089" heatid="9581" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:29.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Viola Jasmine" gender="F" lastname="Provost" nation="GER" license="329228" athleteid="7045">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.92" entrycourse="SCM" eventid="2089" heatid="9585" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:28.12" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Roman" gender="M" lastname="Roelen" nation="GER" license="283816" athleteid="7047">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.64" entrycourse="SCM" eventid="1749" heatid="9362" lane="2">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:05.64" />
                </ENTRY>
                <ENTRY entrytime="00:18:13.66" eventid="1792" heatid="9406" lane="2" />
                <ENTRY entrytime="00:00:25.31" entrycourse="SCM" eventid="1834" heatid="9450" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:25.31" />
                </ENTRY>
                <ENTRY entrytime="00:09:27.26" eventid="2168" status="RJC" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Luis" gender="M" lastname="Steinmassl" nation="GER" license="201458" athleteid="7052">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.05" entrycourse="SCM" eventid="1749" heatid="9364" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:51.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.97" entrycourse="SCM" eventid="1778" heatid="9392" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:54.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.20" entrycourse="SCM" eventid="1834" heatid="9452" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-01-13" name="34. Augsburger Zirbelnuss-Schwimmen" qualificationtime="00:00:23.37" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.25" entrycourse="SCM" eventid="1971" heatid="9495" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-01-12" name="34. Augsburger Zirbelnuss-Schwimmen" qualificationtime="00:00:51.64" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.20" entrycourse="SCM" eventid="2041" heatid="9558" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:07.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.30" entrycourse="SCM" eventid="5307" heatid="9599" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:25.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Steven" gender="M" lastname="Stöckl" nation="GER" license="316820" athleteid="7059">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.69" entrycourse="SCM" eventid="1749" heatid="9365" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:02.69" />
                </ENTRY>
                <ENTRY entrytime="00:17:42.22" entrycourse="SCM" eventid="1792" heatid="9407" lane="1">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:17:42.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.28" entrycourse="SCM" eventid="1834" heatid="9446" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:26.28" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.71" entrycourse="SCM" eventid="1848" heatid="9468" lane="1">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:18.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.64" entrycourse="SCM" eventid="1971" heatid="9491" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:56.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.44" entrycourse="SCM" eventid="2013" heatid="9535" lane="4">
                  <MEETINFO city="Dachau" course="SCM" date="2019-02-10" name="Kreisjahrgangsmeisterschaften Kreis4 Obb." qualificationtime="00:01:03.44" />
                </ENTRY>
                <ENTRY entrytime="00:04:17.67" entrycourse="SCM" eventid="2103" heatid="9612" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:04:17.67" />
                </ENTRY>
                <ENTRY entrytime="00:09:18.89" entrycourse="LCM" eventid="2168" heatid="9616" lane="1">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-03-16" name="International Swim Meeting Erlangen" qualificationtime="00:09:18.89" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Simon" gender="M" lastname="Ulich" nation="GER" license="346570" athleteid="7068">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.20" entrycourse="SCM" eventid="1763" heatid="9383" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:08.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.42" entrycourse="SCM" eventid="1778" heatid="9391" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:01.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.27" entrycourse="SCM" eventid="1985" heatid="9514" lane="1">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:31.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.80" entrycourse="SCM" eventid="2082" heatid="9571" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:26.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.17" entrycourse="SCM" eventid="5307" heatid="9593" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:28.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Antonia" gender="F" lastname="Zerbs" nation="GER" license="351449" athleteid="7074">
              <ENTRIES>
                <ENTRY entrytime="00:20:08.70" entrycourse="LCM" eventid="5318" heatid="9478" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:20:08.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.76" entrycourse="SCM" eventid="1978" heatid="9500" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:20.76" />
                </ENTRY>
                <ENTRY entrytime="00:10:30.34" entrycourse="LCM" eventid="2020" heatid="9541" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-11" name="Erlanger Sparkassen-Cup" qualificationtime="00:10:30.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.63" eventid="5316" heatid="9480" lane="4" />
                <ENTRY entrytime="00:01:45.63" eventid="2232" heatid="9619" lane="2" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.59" eventid="5314" heatid="9482" lane="2" />
                <ENTRY entrytime="00:01:56.33" eventid="2224" heatid="9618" lane="6" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.76" eventid="1855" heatid="9477" lane="6">
                  <MEETINFO city="Kaufering" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:00.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.11" eventid="5303" heatid="9615" lane="6">
                  <MEETINFO city="Kaufering" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:07.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.27" eventid="1855" heatid="9476" lane="4">
                  <MEETINFO city="Kaufering" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:00.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.55" eventid="5303" heatid="9614" lane="5">
                  <MEETINFO city="Kaufering" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:07.91" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6777" nation="GER" region="02" clubid="5735" name="Schwimmclub Schwandorf">
          <CONTACT city="Schwandorf" email="tobias.schwendner@schwimmclub-schwandorf.de" name="Schwendner, Tobias" phone="09431-5283551" street="Föhrenstraße 5" zip="92421" />
          <ATHLETES>
            <ATHLETE birthdate="2001-01-01" firstname="Anika" gender="F" lastname="Jacksteit" nation="GER" license="266125" athleteid="5736">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.39" entrycourse="SCM" eventid="2034" heatid="9553" lane="6">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:00:32.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.86" entrycourse="SCM" eventid="2089" heatid="9583" lane="6">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:00:28.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4302" nation="GER" region="02" clubid="5671" name="Schwimmfreunde Pegnitz">
          <ATHLETES>
            <ATHLETE birthdate="1995-01-01" firstname="Sandra" gender="F" lastname="Bauer" nation="GER" license="197004" athleteid="5672">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.40" entrycourse="SCM" eventid="1756" heatid="9373" lane="4">
                  <MEETINFO city="Pegnitz" course="SCM" date="2019-10-05" name="2. CabrioSol Cup" qualificationtime="00:00:34.40" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.63" entrycourse="SCM" eventid="1799" heatid="9412" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:10.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6399" nation="GER" region="02" clubid="6478" name="SG - Elsenfeld/Kleinwallstadt">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Adriana" gender="F" lastname="Bethke" nation="GER" license="307751" athleteid="6479">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.94" entrycourse="SCM" eventid="2089" heatid="9578" lane="6">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-07-21" name="Kinder- und Jugendschwimmfest" qualificationtime="00:00:29.94" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5085" nation="GER" region="02" clubid="6696" name="SG Bamberg">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Nikita" gender="F" lastname="Bergmann" nation="GER" license="335717" athleteid="6697">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.66" entrycourse="SCM" eventid="1756" heatid="9374" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:34.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.30" entrycourse="SCM" eventid="1827" heatid="9439" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:43.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.73" entrycourse="SCM" eventid="1992" heatid="9522" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:13.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.90" entrycourse="SCM" eventid="2089" heatid="9578" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:29.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Leila" gender="F" lastname="Jafoui" nation="GER" license="342435" athleteid="6702">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.46" entrycourse="SCM" eventid="1756" heatid="9370" lane="4">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-16" name="10. Internationales Frühjahresmeeting" qualificationtime="00:00:36.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.77" entrycourse="SCM" eventid="1799" heatid="9409" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:13.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.86" entrycourse="SCM" eventid="1827" heatid="9436" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:55.86" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.95" entrycourse="SCM" eventid="1992" heatid="9520" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:19.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Kevin" gender="M" lastname="Kertész" nation="GER" license="391557" athleteid="6707">
              <ENTRIES>
                <ENTRY entrytime="00:02:14.61" entrycourse="SCM" eventid="1848" heatid="9467" lane="4">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:02:14.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.55" entrycourse="SCM" eventid="2013" heatid="9537" lane="1">
                  <MEETINFO city="Wetzlar" course="LCM" date="2019-05-04" name="27. Süddeutsche Jahrgangsmeisterschaften" qualificationtime="00:01:03.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Josefin" gender="F" lastname="Krefft" nation="GER" license="361625" athleteid="6710">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.65" entrycourse="SCM" eventid="1059" heatid="9347" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:03.65" />
                </ENTRY>
                <ENTRY entrytime="00:04:56.46" entrycourse="SCM" eventid="5320" heatid="9472" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:04:56.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.69" entrycourse="SCM" eventid="1978" heatid="9501" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:20.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.95" entrycourse="SCM" eventid="2089" heatid="9582" lane="1">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:28.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Maja" gender="F" lastname="Lehner" nation="GER" license="290695" athleteid="6715">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.02" entrycourse="SCM" eventid="1059" heatid="9350" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:02.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.69" entrycourse="SCM" eventid="2006" heatid="9530" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:08.69" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Isabel" gender="F" lastname="Linß" nation="GER" license="165184" athleteid="6718">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.14" entrycourse="SCM" eventid="1799" heatid="9411" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:11.14" />
                </ENTRY>
                <ENTRY entrytime="00:04:48.86" entrycourse="SCM" eventid="5320" heatid="9473" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:04:48.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.26" entrycourse="SCM" eventid="1978" heatid="9503" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:16.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.66" entrycourse="SCM" eventid="1992" heatid="9523" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:17.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.87" entrycourse="SCM" eventid="2089" heatid="9582" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:28.87" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Bastian" gender="M" lastname="Schorr" nation="GER" license="137664" athleteid="6724">
              <ENTRIES>
                <ENTRY entrytime="00:01:55.00" entrycourse="SCM" eventid="1749" heatid="9363" lane="4">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:01:52.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.50" entrycourse="SCM" eventid="1834" heatid="9454" lane="6">
                  <MEETINFO city="Pegnitz" course="SCM" date="2019-10-05" name="2. CabrioSol Cup" qualificationtime="00:00:24.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.00" entrycourse="SCM" eventid="1971" heatid="9494" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:00:54.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.00" entrycourse="SCM" eventid="5307" heatid="9598" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:00:26.49" />
                </ENTRY>
                <ENTRY entrytime="00:04:15.00" entrycourse="SCM" eventid="2103" heatid="9613" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:04:17.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Gregor" gender="M" lastname="Spörlein" nation="GER" license="158773" athleteid="6730">
              <ENTRIES>
                <ENTRY entrytime="00:01:48.70" entrycourse="SCM" eventid="1749" heatid="9365" lane="3">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:01:48.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.09" entrycourse="SCM" eventid="1778" heatid="9393" lane="3">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:00:54.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.74" entrycourse="SCM" eventid="1834" heatid="9452" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-04" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:00:23.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.32" entrycourse="SCM" eventid="1971" heatid="9497" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-04" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:00:51.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.64" entrycourse="SCM" eventid="2041" heatid="9559" lane="3">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:02:03.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.01" entrycourse="SCM" eventid="5307" heatid="9598" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-04" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:00:25.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Martin" gender="M" lastname="Spörlein" nation="GER" license="169787" athleteid="6737">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.79" entrycourse="SCM" eventid="1749" heatid="9365" lane="1">
                  <MEETINFO city="Essen" course="LCM" date="2019-05-11" name="German Open im Schwimmen" qualificationtime="00:02:00.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.60" entrycourse="SCM" eventid="1834" heatid="9454" lane="3">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:00:22.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.45" entrycourse="SCM" eventid="1971" heatid="9496" lane="4">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:00:51.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.34" entrycourse="SCM" eventid="5307" heatid="9595" lane="6">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:27.34" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Ella" gender="F" lastname="Vornlocher" nation="GER" license="335716" athleteid="6742">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.05" entrycourse="SCM" eventid="2089" heatid="9576" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:30.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.10" eventid="5316" heatid="9481" lane="5">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:55.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.70" eventid="2232" heatid="9620" lane="4">
                  <MEETINFO city="Kulmbach" date="2019-02-16" name="6. Kulmbacher-Kinder-Schwimm-Vergnügen" qualificationtime="00:03:06.98" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.80" eventid="1855" heatid="9477" lane="5">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:49.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:58.80" eventid="5303" heatid="9614" lane="3">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:02:02.94" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5068" nation="GER" region="02" clubid="5815" name="SG Haßberge">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Johanna" gender="F" lastname="Strobel" nation="GER" license="334239" athleteid="5816">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.26" entrycourse="SCM" eventid="1799" heatid="9408" lane="3">
                  <MEETINFO city="Lohr am Main" course="SCM" date="2019-03-23" name="Ufr.- &amp; 2. intern. Master-Kurzbahnmeisterschaften" qualificationtime="00:01:14.77" />
                </ENTRY>
                <ENTRY entrytime="00:02:50.64" entrycourse="SCM" eventid="1827" heatid="9438" lane="1">
                  <MEETINFO city="Haßfurt" course="SCM" date="2019-02-03" name="Kreismeisterschaft Kreis Main-Rhön  Kurzbahn" qualificationtime="00:02:50.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.21" entrycourse="SCM" eventid="1992" heatid="9521" lane="1">
                  <MEETINFO city="Schweinfurt" course="SCM" date="2019-01-19" name="10. Juki Schwimmfest" qualificationtime="00:01:19.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5212" nation="GER" region="02" clubid="5675" name="SG Mallersdorf/Pfaffenberg">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Christina" gender="F" lastname="Gockeln" nation="GER" license="342662" athleteid="5676">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.18" entrycourse="SCM" eventid="1992" heatid="9521" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-31" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:01:19.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julian" gender="M" lastname="Gockeln" nation="GER" license="342661" athleteid="5678">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.48" entrycourse="SCM" eventid="1985" heatid="9512" lane="5">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:32.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Simon" gender="M" lastname="Koci" nation="GER" license="353012" athleteid="5680">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.63" entrycourse="SCM" eventid="1971" heatid="9489" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-03-30" name="Ndb. Kurzbahnmeisterschaften Jahrg. 2011 u. ällter" qualificationtime="00:00:57.63" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.31" entrycourse="SCM" eventid="5307" heatid="9593" lane="2">
                  <MEETINFO city="Neustadt/Donau" course="SCM" date="2019-03-17" name="Ndb. Kreismeisterschaften West" qualificationtime="00:00:28.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6768" nation="GER" region="02" clubid="6752" name="SG Mittelfranken">
          <ATHLETES>
            <ATHLETE birthdate="2006-01-01" firstname="Michael" gender="M" lastname="Bachmann" nation="GER" license="354895" athleteid="6753">
              <ENTRIES>
                <ENTRY entrytime="00:04:37.10" entrycourse="LCM" eventid="2103" heatid="9609" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:44.31" />
                </ENTRY>
                <ENTRY entrytime="00:09:35.83" entrycourse="LCM" eventid="2168" heatid="9616" lane="6">
                  <MEETINFO city="Kleinostheim" course="LCM" date="2019-05-04" name="Nationales Schwimm-Meeting" qualificationtime="00:09:50.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Anna" gender="F" lastname="Baumgarte" nation="GER" license="331994" athleteid="6756">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.75" entrycourse="SCM" eventid="1059" heatid="9346" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:05.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.63" entrycourse="SCM" eventid="1978" heatid="9502" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:20.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.43" entrycourse="SCM" eventid="2089" heatid="9579" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:29.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Lorenz" gender="M" lastname="Beck" nation="GER" license="337791" athleteid="6760">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.99" entrycourse="SCM" eventid="1763" heatid="9379" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-01-26" name="DSV Endkampf DMSJ" qualificationtime="00:01:12.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.63" entrycourse="SCM" eventid="1778" heatid="9390" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:02.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.60" entrycourse="SCM" eventid="1820" heatid="9433" lane="6">
                  <MEETINFO city="Wetzlar" course="LCM" date="2019-05-04" name="27. Süddeutsche Jahrgangsmeisterschaften" qualificationtime="00:02:23.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.97" entrycourse="SCM" eventid="1985" heatid="9511" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:32.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.51" entrycourse="SCM" eventid="2027" heatid="9545" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:04.51" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.65" entrycourse="SCM" eventid="2082" heatid="9570" lane="4">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:35.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Reka" gender="F" lastname="Behring" nation="GER" license="313608" athleteid="6767">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.14" entrycourse="SCM" eventid="2034" heatid="9555" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:32.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.35" entrycourse="SCM" eventid="2089" heatid="9587" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:27.35" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.76" entrycourse="SCM" eventid="2096" heatid="9604" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:32.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Thomas" gender="M" lastname="Chang" nation="GER" license="201143" athleteid="6771">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.29" entrycourse="SCM" eventid="1763" heatid="9381" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:09.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.38" entrycourse="SCM" eventid="1971" heatid="9491" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:56.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lisa" gender="F" lastname="Emmerlich-Mace" nation="GER" license="390428" athleteid="6774">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.83" entrycourse="SCM" eventid="1785" heatid="9398" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:12.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.63" entrycourse="SCM" eventid="2034" heatid="9550" lane="3">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:33.63" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.84" entrycourse="SCM" eventid="2096" heatid="9603" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:34.84" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Taliso" gender="M" lastname="Engel" nation="GER" license="282421" athleteid="6778">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.25" entrycourse="SCM" eventid="1763" heatid="9382" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:06.25" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.14" entrycourse="SCM" eventid="1820" heatid="9433" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:02:21.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.12" entrycourse="LCM" eventid="1834" heatid="9447" lane="2">
                  <MEETINFO city="Hannover" course="LCM" date="2019-02-23" name="21. Piranha-Meeting" qualificationtime="00:00:26.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.70" entrycourse="LCM" eventid="1971" heatid="9490" lane="3">
                  <MEETINFO city="Hannover" course="LCM" date="2019-02-24" name="21. Piranha-Meeting" qualificationtime="00:00:58.52" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.31" entrycourse="LCM" eventid="1985" heatid="9516" lane="4">
                  <MEETINFO city="Hannover" course="LCM" date="2019-02-24" name="21. Piranha-Meeting" qualificationtime="00:00:30.31" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.62" entrycourse="SCM" eventid="2082" heatid="9573" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:02:27.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.00" eventid="5307" heatid="9596" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sofia Lucia" gender="F" lastname="Giurbino" nation="GER" license="319882" athleteid="6786">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.88" entrycourse="SCM" eventid="1059" heatid="9345" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:05.88" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.53" entrycourse="SCM" eventid="1756" heatid="9370" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:36.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.03" entrycourse="SCM" eventid="2089" heatid="9577" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:30.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1993-01-01" firstname="Daniela" gender="F" lastname="Karst" nation="GER" license="156320" athleteid="6790">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.00" entrycourse="SCM" eventid="1756" heatid="9374" lane="3">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:33.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.50" entrycourse="SCM" eventid="1799" heatid="9414" lane="3">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:10.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.50" entrycourse="SCM" eventid="1841" heatid="9463" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-05-25" name="Deutsche Hochschulmeisterschaften" qualificationtime="00:00:28.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.00" entrycourse="SCM" eventid="2006" heatid="9530" lane="3">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:01:02.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.90" entrycourse="SCM" eventid="2089" heatid="9587" lane="3">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:00:27.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Clemens" gender="M" lastname="Knorr" nation="GER" license="326926" athleteid="6796">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.39" entrycourse="SCM" eventid="1971" heatid="9485" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:59.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Oliver" gender="M" lastname="Kreißel" nation="GER" license="313677" athleteid="6801">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.56" entrycourse="SCM" eventid="1763" heatid="9384" lane="6">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:09.51" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.87" entrycourse="SCM" eventid="1778" heatid="9391" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:02.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.47" entrycourse="SCM" eventid="1820" heatid="9432" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:17.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.18" entrycourse="SCM" eventid="1971" heatid="9485" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:00:59.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.80" entrycourse="SCM" eventid="1985" heatid="9516" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:30.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.91" entrycourse="SCM" eventid="2027" heatid="9546" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:02.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.83" entrycourse="LCM" eventid="2082" heatid="9573" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:38.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Ira" gender="F" lastname="Ködel" nation="GER" license="295234" athleteid="6798">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.00" entrycourse="SCM" eventid="1785" heatid="9397" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:14.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Michelle" gender="F" lastname="Messel" nation="GER" license="196996" athleteid="6809">
              <ENTRIES>
                <ENTRY entrytime="00:02:28.00" entrycourse="SCM" eventid="1813" heatid="9425" lane="2">
                  <MEETINFO city="Amberg" course="LCM" date="2019-06-02" name="Kurfürstenpokal" qualificationtime="00:02:24.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.50" entrycourse="SCM" eventid="1841" heatid="9463" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:29.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.50" entrycourse="SCM" eventid="2006" heatid="9531" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:05.97" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.80" entrycourse="SCM" eventid="2034" heatid="9552" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:31.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Marvin" gender="M" lastname="Metz" nation="GER" license="323026" athleteid="6814">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.90" entrycourse="SCM" eventid="1749" heatid="9359" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:02:07.90" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.03" entrycourse="SCM" eventid="1834" heatid="9447" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:00:26.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.28" entrycourse="SCM" eventid="1971" heatid="9487" lane="4">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:58.09" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.59" entrycourse="SCM" eventid="2013" heatid="9534" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Ingolstadt" qualificationtime="00:01:06.59" />
                </ENTRY>
                <ENTRY entrytime="00:04:30.74" entrycourse="LCM" eventid="2103" heatid="9610" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:30.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Luna" gender="F" lastname="Ohlschmid" nation="GER" license="331164" athleteid="6820">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.70" entrycourse="SCM" eventid="1756" heatid="9371" lane="3">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:37.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Jeremias" gender="M" lastname="Pock" nation="GER" license="269306" athleteid="6822">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.81" entrycourse="SCM" eventid="1763" heatid="9384" lane="4">
                  <MEETINFO city="Mainz" course="SCM" date="2019-02-02" name="DMS 2. Bundesliga Süd" qualificationtime="00:01:06.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.78" entrycourse="LCM" eventid="1778" heatid="9394" lane="4">
                  <MEETINFO city="Nürnberg" course="LCM" date="2019-07-06" name="Mittelfränkische Meisterschaften" qualificationtime="00:00:59.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.31" entrycourse="SCM" eventid="1820" heatid="9432" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:08.31" />
                </ENTRY>
                <ENTRY entrytime="00:04:38.87" entrycourse="SCM" eventid="1999" heatid="9527" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:04:40.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.10" entrycourse="SCM" eventid="2027" heatid="9546" lane="3">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:59.42" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.75" entrycourse="SCM" eventid="2082" heatid="9571" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:22.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.70" entrycourse="SCM" eventid="5307" heatid="9597" lane="4">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:26.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Laura" gender="F" lastname="Popp" nation="GER" license="178550" athleteid="6830">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.00" entrycourse="SCM" eventid="1992" heatid="9523" lane="4">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:16.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:32.00" entrycourse="LCM" eventid="2075" heatid="9565" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-11" name="Erlanger Sparkassen-Cup" qualificationtime="00:02:34.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Charlotte" gender="F" lastname="Rudat" nation="GER" license="330018" athleteid="6833">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.22" entrycourse="SCM" eventid="1841" heatid="9462" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:30.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.91" entrycourse="SCM" eventid="2034" heatid="9552" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:32.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.95" entrycourse="SCM" eventid="2089" heatid="9585" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:27.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Jan" gender="M" lastname="Sedlacek" nation="GER" license="315494" athleteid="6865">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.90" entrycourse="SCM" eventid="1763" heatid="9377" lane="1">
                  <MEETINFO city="Frankenberg (Eder)" course="SCM" date="2019-05-04" name="49. Int. Maischwimmen" qualificationtime="00:01:14.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.80" entrycourse="SCM" eventid="1820" heatid="9429" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:25.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.30" entrycourse="SCM" eventid="1985" heatid="9509" lane="1">
                  <MEETINFO city="Forchheim" course="SCM" date="2019-03-23" name="16. Frühjahrs-Sprint-Meeting_Ausschreibung" qualificationtime="00:00:33.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:42.10" entrycourse="SCM" eventid="2082" heatid="9570" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:41.67" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Nele" gender="F" lastname="Sturm" nation="GER" license="297331" athleteid="6837">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.15" entrycourse="LCM" eventid="1756" heatid="9372" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:34.18" />
                </ENTRY>
                <ENTRY entrytime="00:05:14.05" entrycourse="LCM" eventid="1771" heatid="9388" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:05:14.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.24" entrycourse="LCM" eventid="1827" heatid="9437" lane="2">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:02:47.54" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.82" entrycourse="SCM" eventid="1992" heatid="9523" lane="2">
                  <MEETINFO city="Essen" course="SCM" date="2019-01-26" name="DSV Endkampf DMSJ" qualificationtime="00:01:15.82" />
                </ENTRY>
                <ENTRY entrytime="00:09:37.23" entrycourse="LCM" eventid="2020" heatid="9541" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:09:37.23" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.44" entrycourse="LCM" eventid="2075" heatid="9566" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:31.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lucy" gender="F" lastname="Suljewic" nation="GER" license="316692" athleteid="6844">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.99" entrycourse="SCM" eventid="1059" heatid="9348" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:02.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.62" entrycourse="SCM" eventid="1785" heatid="9400" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:10.94" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.37" entrycourse="SCM" eventid="1799" heatid="9410" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:13.31" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.53" entrycourse="SCM" eventid="1978" heatid="9502" lane="5">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-12" name="Int. arena Swim Meeting" qualificationtime="00:02:18.68" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.17" entrycourse="SCM" eventid="2034" heatid="9553" lane="1">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:33.06" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.17" entrycourse="SCM" eventid="2089" heatid="9581" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:29.17" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.60" entrycourse="SCM" eventid="2096" heatid="9606" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:29.80" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Julian" gender="M" lastname="Vogl" nation="GER" license="358408" athleteid="6852">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.50" entrycourse="SCM" eventid="1763" heatid="9380" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:10.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.89" entrycourse="SCM" eventid="1834" heatid="9448" lane="3">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:25.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.43" entrycourse="SCM" eventid="1971" heatid="9489" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:57.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.92" entrycourse="SCM" eventid="1985" heatid="9515" lane="5">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:30.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Rebecca" gender="F" lastname="Walther" nation="GER" license="292203" athleteid="6857">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.30" entrycourse="SCM" eventid="1756" heatid="9373" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:35.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:18.37" entrycourse="SCM" eventid="1992" heatid="9521" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:18.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Marie" gender="F" lastname="Wormser" nation="GER" license="292535" athleteid="6860">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.71" entrycourse="SCM" eventid="1799" heatid="9411" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:11.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.26" entrycourse="SCM" eventid="2034" heatid="9554" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:32.26" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Natalie" gender="F" lastname="Wöltinger" nation="GER" license="266843" athleteid="6890">
              <ENTRIES>
                <ENTRY entrytime="00:04:59.90" entrycourse="SCM" eventid="1771" heatid="9388" lane="4">
                  <MEETINFO city="Wiesbaden" course="SCM" date="2019-02-02" name="DMS Oberliga Hessen" qualificationtime="00:04:59.90" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.05" entrycourse="LCM" eventid="1827" heatid="9437" lane="3">
                  <MEETINFO city="Kassel" course="LCM" date="2019-06-01" name="35.Schwimmfest" qualificationtime="00:02:47.11" />
                </ENTRY>
                <ENTRY entrytime="00:04:25.67" entrycourse="LCM" eventid="5320" heatid="9475" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-02" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:04:34.81" />
                </ENTRY>
                <ENTRY entrytime="00:09:39.54" entrycourse="LCM" eventid="2020" heatid="9541" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-02-24" name="30. Süddeutsche Meisterschaften Lange Strecken" qualificationtime="00:09:39.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.41" entrycourse="SCM" eventid="2075" heatid="9565" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-03" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:02:24.09" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.19" eventid="2232" heatid="9620" lane="3" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:46.27" eventid="5303" heatid="9615" lane="3" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="5541" nation="GER" region="02" clubid="5844" name="SG Nordoberpfalz">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Kathrin" gender="F" lastname="Bachmeier" nation="GER" license="262269" athleteid="5845">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.82" entrycourse="SCM" eventid="1059" heatid="9355" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:59.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.58" entrycourse="SCM" eventid="1799" heatid="9414" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:09.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.62" entrycourse="SCM" eventid="1841" heatid="9462" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:29.62" />
                </ENTRY>
                <ENTRY entrytime="00:04:35.60" entrycourse="SCM" eventid="5320" heatid="9475" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:46.46" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.56" entrycourse="SCM" eventid="1978" heatid="9506" lane="4">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:11.08" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.20" entrycourse="SCM" eventid="2006" heatid="9530" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:07.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.26" entrycourse="SCM" eventid="2089" heatid="9588" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:27.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Viktoria" gender="F" lastname="Bogner" nation="GER" license="287903" athleteid="5853">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.73" entrycourse="SCM" eventid="1059" heatid="9355" lane="1">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:59.73" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.00" entrycourse="SCM" eventid="1799" heatid="9411" lane="3">
                  <MEETINFO city="Plauen" course="SCM" date="2019-09-28" name="Plauener Herbst-Mehrkampf" qualificationtime="00:01:11.00" />
                </ENTRY>
                <ENTRY entrytime="00:04:46.38" entrycourse="SCM" eventid="5320" heatid="9474" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:04:48.61" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.11" entrycourse="SCM" eventid="1978" heatid="9505" lane="2">
                  <MEETINFO city="Tirschenreuth" course="SCM" date="2019-04-28" name="17. Internationale Frühlingsschwimmen mit kindgere" qualificationtime="00:02:11.11" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.57" entrycourse="SCM" eventid="2075" heatid="9567" lane="6">
                  <MEETINFO city="Tirschenreuth" course="SCM" date="2019-04-28" name="17. Internationale Frühlingsschwimmen mit kindgere" qualificationtime="00:02:31.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.82" entrycourse="SCM" eventid="2089" heatid="9586" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:27.90" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Daria" gender="F" lastname="Codlova" nation="GER" license="356592" athleteid="5860">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.15" entrycourse="SCM" eventid="1756" heatid="9369" lane="2">
                  <MEETINFO city="Tirschenreuth" course="SCM" date="2019-04-28" name="17. Internationale Frühlingsschwimmen mit kindgere" qualificationtime="00:00:37.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Fynn" gender="M" lastname="Legat" nation="GER" license="339495" athleteid="5862">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.03" entrycourse="SCM" eventid="1763" heatid="9378" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:13.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.48" entrycourse="SCM" eventid="1985" heatid="9512" lane="2">
                  <MEETINFO city="Tirschenreuth" course="SCM" date="2019-04-28" name="17. Internationale Frühlingsschwimmen mit kindgere" qualificationtime="00:00:32.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Kilian" gender="M" lastname="Züllich" nation="GER" license="262780" athleteid="5865">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.36" entrycourse="SCM" eventid="1763" heatid="9379" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:12.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.08" entrycourse="SCM" eventid="1985" heatid="9513" lane="2">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:32.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4305" nation="GER" region="02" clubid="6481" name="SG Oberland Penzberg">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Nele" gender="F" lastname="Bäck" nation="GER" license="318082" athleteid="6482">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.50" entrycourse="SCM" eventid="1756" heatid="9368" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:37.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sara" gender="F" lastname="Lickel" nation="GER" license="322797" athleteid="6484">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.57" entrycourse="SCM" eventid="2034" heatid="9551" lane="1">
                  <MEETINFO city="Kaufbeuren" course="SCM" date="2019-03-24" name="18. Internationaler Buron Cup" qualificationtime="00:00:33.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6423" nation="GER" region="02" clubid="6055" name="SG Stadtwerke München">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Ivan" gender="M" lastname="Anzarski" nation="GER" license="368146" athleteid="6056">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.04" entrycourse="SCM" eventid="1763" heatid="9383" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:07.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.85" entrycourse="SCM" eventid="1820" heatid="9431" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:17.85" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.84" entrycourse="SCM" eventid="1971" heatid="9490" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:56.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.97" entrycourse="SCM" eventid="1985" heatid="9514" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:30.97" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.53" eventid="2027" heatid="9544" lane="6" />
                <ENTRY entrytime="00:02:29.48" entrycourse="SCM" eventid="2082" heatid="9572" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:29.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Silvian" gender="M" lastname="Balbach" nation="GER" license="315759" athleteid="6063">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.64" entrycourse="SCM" eventid="1749" heatid="9363" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:02.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.91" entrycourse="SCM" eventid="1778" heatid="9389" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:02.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.74" entrycourse="SCM" eventid="1820" heatid="9432" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:21.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.94" entrycourse="SCM" eventid="1834" heatid="9451" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:24.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.81" entrycourse="SCM" eventid="1971" heatid="9492" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:55.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.29" eventid="2027" heatid="9543" lane="1" />
                <ENTRY entrytime="00:00:28.35" entrycourse="SCM" eventid="5307" heatid="9593" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:28.35" />
                </ENTRY>
                <ENTRY entrytime="00:04:24.57" entrycourse="SCM" eventid="2103" heatid="9612" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:04:24.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Yael" gender="M" lastname="Balz" nation="GER" license="318639" athleteid="6072">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.53" entrycourse="LCM" eventid="1749" heatid="9364" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:59.27" />
                </ENTRY>
                <ENTRY entrytime="00:16:26.35" entrycourse="SCM" eventid="1792" heatid="9407" lane="4">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:16:39.30" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.09" entrycourse="SCM" eventid="1820" heatid="9432" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:16.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.90" entrycourse="SCM" eventid="1971" heatid="9496" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:55.60" />
                </ENTRY>
                <ENTRY entrytime="00:04:05.89" entrycourse="LCM" eventid="2103" heatid="9613" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:13.47" />
                </ENTRY>
                <ENTRY entrytime="00:08:32.45" entrycourse="LCM" eventid="2168" heatid="9617" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-15" name="10. Internationales Frühjahresmeeting" qualificationtime="00:08:51.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1973-01-01" firstname="Markus" gender="M" lastname="Bierig" nation="GER" license="56866" athleteid="6079">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" entrycourse="SCM" eventid="1778" heatid="9393" lane="1">
                  <MEETINFO city="Karlsruhe" course="LCM" date="2019-06-01" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:01:00.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.00" entrycourse="SCM" eventid="1971" heatid="9492" lane="2">
                  <MEETINFO city="Dachau" course="SCM" date="2019-02-16" name="20. Int. Dachauer Masters-Cup" qualificationtime="00:00:56.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.50" entrycourse="SCM" eventid="5307" heatid="9598" lane="1">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:26.60" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Moritz" gender="M" lastname="Bockes" nation="GER" license="279879" athleteid="6083">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.99" entrycourse="SCM" eventid="1749" heatid="9364" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:03.96" />
                </ENTRY>
                <ENTRY entrytime="00:16:43.40" entrycourse="SCM" eventid="1792" heatid="9407" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:16:43.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.25" entrycourse="SCM" eventid="1971" heatid="9489" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:57.25" />
                </ENTRY>
                <ENTRY entrytime="00:04:15.92" entrycourse="SCM" eventid="2103" heatid="9612" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:15.92" />
                </ENTRY>
                <ENTRY entrytime="00:08:52.52" entrycourse="LCM" eventid="2168" heatid="9617" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:08:52.52" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Pascal" gender="M" lastname="Borchardt" nation="GER" license="287497" athleteid="6089">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.00" entrycourse="SCM" eventid="1778" heatid="9393" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:00.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.45" entrycourse="SCM" eventid="1806" heatid="9420" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:27.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.37" eventid="1834" heatid="9453" lane="5" />
                <ENTRY entrytime="00:00:52.79" entrycourse="SCM" eventid="1971" heatid="9495" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:55.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.46" eventid="2013" heatid="9537" lane="4" />
                <ENTRY entrytime="00:01:00.54" eventid="2027" heatid="9546" lane="4" />
                <ENTRY entrytime="00:00:26.46" eventid="5307" heatid="9597" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Manuel" gender="M" lastname="Cubero" nation="GER" license="353771" athleteid="6097">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.74" entrycourse="SCM" eventid="1834" heatid="9452" lane="6">
                  <MEETINFO city="Dortmund" course="LCM" date="2019-03-16" name="20. Internationales Sparkassen ISDO" qualificationtime="00:00:24.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.07" entrycourse="SCM" eventid="1971" heatid="9490" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:57.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.47" entrycourse="LCM" eventid="5307" heatid="9593" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-12" name="Erlanger Sparkassen-Cup" qualificationtime="00:00:28.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Henning" gender="M" lastname="Dörries" nation="GER" license="220261" athleteid="6101">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.12" entrycourse="LCM" eventid="1749" heatid="9365" lane="4">
                  <MEETINFO city="Merano" course="LCM" date="2019-06-29" name="Cool Swim Meeting" qualificationtime="00:01:59.42" />
                </ENTRY>
                <ENTRY entrytime="00:15:55.00" entrycourse="SCM" eventid="1792" heatid="9407" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:16:04.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.84" entrycourse="SCM" eventid="1820" heatid="9431" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:13.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.86" entrycourse="SCM" eventid="1971" heatid="9497" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:54.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.49" eventid="2041" heatid="9558" lane="5" />
                <ENTRY entrytime="00:02:17.79" entrycourse="SCM" eventid="2082" heatid="9573" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-03" name="DMS 1. Bundesliga" qualificationtime="00:02:19.97" />
                </ENTRY>
                <ENTRY entrytime="00:04:00.23" entrycourse="SCM" eventid="2103" heatid="9613" lane="4">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:04:03.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Luise" gender="F" lastname="Dörries" nation="GER" license="162166" athleteid="6109">
              <ENTRIES>
                <ENTRY entrytime="00:02:24.45" entrycourse="LCM" eventid="1813" heatid="9425" lane="4">
                  <MEETINFO city="Merano" course="LCM" date="2019-06-28" name="Cool Swim Meeting" qualificationtime="00:02:28.08" />
                </ENTRY>
                <ENTRY entrytime="00:04:34.87" entrycourse="LCM" eventid="5320" heatid="9475" lane="5">
                  <MEETINFO city="Merano" course="LCM" date="2019-06-28" name="Cool Swim Meeting" qualificationtime="00:04:37.62" />
                </ENTRY>
                <ENTRY entrytime="00:17:12.20" entrycourse="LCM" eventid="5318" heatid="9479" lane="3">
                  <MEETINFO city="Merano" course="LCM" date="2019-06-29" name="Cool Swim Meeting" qualificationtime="00:17:39.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.74" entrycourse="LCM" eventid="1978" heatid="9506" lane="6">
                  <MEETINFO city="Merano" course="LCM" date="2019-06-29" name="Cool Swim Meeting" qualificationtime="00:02:15.47" />
                </ENTRY>
                <ENTRY entrytime="00:09:08.01" entrycourse="LCM" eventid="2020" heatid="9541" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:09:20.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Manuel" gender="M" lastname="Genster" nation="GER" license="240652" athleteid="6123">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.14" eventid="1749" heatid="9364" lane="4" />
                <ENTRY entrytime="00:00:53.68" entrycourse="SCM" eventid="1778" heatid="9394" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-01" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:00:55.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.93" entrycourse="SCM" eventid="1834" heatid="9453" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:00:22.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:50.42" entrycourse="SCM" eventid="1971" heatid="9497" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:00:50.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.39" entrycourse="LCM" eventid="5307" heatid="9599" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-04" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:00:25.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Rabea" gender="F" lastname="Gärtner" nation="GER" license="316345" athleteid="6115">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.83" entrycourse="LCM" eventid="1059" heatid="9349" lane="1">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:01:02.83" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.00" eventid="1799" heatid="9414" lane="2" />
                <ENTRY entrytime="00:00:30.94" entrycourse="LCM" eventid="1841" heatid="9458" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:30.94" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.23" entrycourse="LCM" eventid="1978" heatid="9501" lane="4">
                  <MEETINFO city="Dortmund" course="LCM" date="2019-03-16" name="20. Internationales Sparkassen ISDO" qualificationtime="00:02:19.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.27" entrycourse="LCM" eventid="2006" heatid="9531" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:07.27" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.72" entrycourse="SCM" eventid="2075" heatid="9565" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:29.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.75" entrycourse="LCM" eventid="2096" heatid="9603" lane="3">
                  <MEETINFO city="Graz-Eggenberg" course="LCM" date="2019-04-26" name="Int. Ströck ATUS Graz Trophy" qualificationtime="00:02:34.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Saskia" gender="F" lastname="Hahn" nation="GER" license="223350" athleteid="6129">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.53" entrycourse="SCM" eventid="1059" heatid="9354" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:00.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.96" entrycourse="SCM" eventid="1813" heatid="9425" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-03" name="DMS 1. Bundesliga" qualificationtime="00:02:18.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.53" entrycourse="SCM" eventid="2006" heatid="9531" lane="4">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:01:04.53" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.34" entrycourse="SCM" eventid="2075" heatid="9566" lane="4">
                  <MEETINFO city="Halle (Saale)" course="LCM" date="2019-03-23" name="19. Schwimmfest" qualificationtime="00:02:26.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Mia" gender="F" lastname="Heinrichsdorff" nation="GER" license="376340" athleteid="6134">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.83" entrycourse="SCM" eventid="1059" heatid="9349" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:01:02.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.40" entrycourse="SCM" eventid="1785" heatid="9403" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:10.31" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.86" eventid="1799" heatid="9412" lane="6" />
                <ENTRY entrytime="00:00:31.44" entrycourse="SCM" eventid="1841" heatid="9458" lane="1">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-12" name="Erlanger Sparkassen-Cup" qualificationtime="00:00:31.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.02" entrycourse="SCM" eventid="2034" heatid="9553" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:33.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.44" entrycourse="SCM" eventid="2075" heatid="9564" lane="1">
                  <MEETINFO city="Graz-Eggenberg" course="LCM" date="2019-04-28" name="Int. Ströck ATUS Graz Trophy" qualificationtime="00:02:34.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.97" entrycourse="SCM" eventid="2089" heatid="9582" lane="6">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:28.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.57" entrycourse="SCM" eventid="2096" heatid="9605" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:30.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Andreas" gender="M" lastname="März" nation="GER" license="301258" athleteid="6143">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.30" entrycourse="SCM" eventid="2013" heatid="9538" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-01-27" name="DSV Endkampf DMSJ" qualificationtime="00:00:56.30" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.65" eventid="2027" heatid="9544" lane="4" />
                <ENTRY entrytime="00:02:10.52" entrycourse="LCM" eventid="2041" heatid="9558" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:10.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.66" entrycourse="SCM" eventid="2082" heatid="9572" lane="4">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:02:25.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Mara" gender="F" lastname="Münsch" nation="GER" license="280574" athleteid="6148">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.50" entrycourse="SCM" eventid="1059" heatid="9352" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:01.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.55" eventid="1799" heatid="9412" lane="4" />
                <ENTRY entrytime="00:02:48.51" entrycourse="SCM" eventid="1827" heatid="9439" lane="5">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:02:52.03" />
                </ENTRY>
                <ENTRY entrytime="00:04:33.03" entrycourse="SCM" eventid="5320" heatid="9475" lane="2">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-03" name="DMS 1. Bundesliga" qualificationtime="00:04:33.03" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.07" entrycourse="LCM" eventid="1978" heatid="9504" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:11.07" />
                </ENTRY>
                <ENTRY entrytime="00:09:28.94" entrycourse="SCM" eventid="2020" heatid="9541" lane="4">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:09:30.55" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Aleksandar" gender="M" lastname="Savic" nation="GER" license="292599" athleteid="6155">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.07" entrycourse="SCM" eventid="1778" heatid="9392" lane="4">
                  <MEETINFO city="Essen" course="SCM" date="2019-01-27" name="DSV Endkampf DMSJ" qualificationtime="00:00:58.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.71" entrycourse="SCM" eventid="1834" heatid="9453" lane="4">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:00:23.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.05" entrycourse="SCM" eventid="1971" heatid="9496" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:00:51.41" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.93" entrycourse="LCM" eventid="2041" heatid="9559" lane="5">
                  <MEETINFO city="Erding" course="LCM" date="2019-07-06" name="Oberbayerische Jahrgangsmeisterschaften" qualificationtime="00:02:19.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.10" entrycourse="LCM" eventid="5307" heatid="9597" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:25.10" />
                </ENTRY>
                <ENTRY entrytime="00:03:58.90" entrycourse="SCM" eventid="2103" heatid="9613" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-03" name="DMS 1. Bundesliga" qualificationtime="00:03:58.90" />
                </ENTRY>
                <ENTRY entrytime="00:08:32.91" entrycourse="LCM" eventid="2168" heatid="9617" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:08:33.58" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Julia" gender="F" lastname="Titze" nation="GER" license="272986" athleteid="6163">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.07" entrycourse="SCM" eventid="1059" heatid="9354" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-04" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:00:57.15" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.92" entrycourse="LCM" eventid="1785" heatid="9402" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-16" name="10. Internationales Frühjahresmeeting" qualificationtime="00:01:08.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.97" eventid="1799" heatid="9415" lane="3" />
                <ENTRY entrytime="00:01:11.17" entrycourse="SCM" eventid="1992" heatid="9524" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-03" name="DMS 1. Bundesliga" qualificationtime="00:01:11.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:17.78" entrycourse="SCM" eventid="2075" heatid="9567" lane="3">
                  <MEETINFO city="Essen" course="SCM" date="2019-02-02" name="DMS 1. Bundesliga" qualificationtime="00:02:18.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.91" entrycourse="LCM" eventid="2089" heatid="9588" lane="4">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-16" name="10. Internationales Frühjahresmeeting" qualificationtime="00:00:27.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lea" gender="F" lastname="Winzer" nation="GER" license="316349" athleteid="6170">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.75" entrycourse="SCM" eventid="1059" heatid="9347" lane="5">
                  <MEETINFO city="Graz-Eggenberg" course="LCM" date="2019-04-28" name="Int. Ströck ATUS Graz Trophy" qualificationtime="00:01:03.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.48" entrycourse="SCM" eventid="1785" heatid="9402" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:09.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.42" eventid="1799" heatid="9410" lane="5" />
                <ENTRY entrytime="00:00:31.08" entrycourse="SCM" eventid="1841" heatid="9458" lane="4">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-12" name="Erlanger Sparkassen-Cup" qualificationtime="00:00:31.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.02" entrycourse="SCM" eventid="1978" heatid="9502" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:19.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.99" entrycourse="SCM" eventid="2034" heatid="9551" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:32.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.21" entrycourse="SCM" eventid="2089" heatid="9580" lane="4">
                  <MEETINFO city="Graz-Eggenberg" course="LCM" date="2019-04-27" name="Int. Ströck ATUS Graz Trophy" qualificationtime="00:00:29.21" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.00" entrycourse="SCM" eventid="2096" heatid="9605" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:29.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Cedric Etienne" gender="M" lastname="Wolf" nation="GER" license="319117" athleteid="6179">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.07" entrycourse="LCM" eventid="1749" heatid="9361" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-12" name="Erlanger Sparkassen-Cup" qualificationtime="00:02:06.07" />
                </ENTRY>
                <ENTRY entrytime="00:17:15.00" entrycourse="SCM" eventid="1792" heatid="9407" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:17:15.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.01" entrycourse="SCM" eventid="1806" heatid="9418" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:30.40" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.32" entrycourse="SCM" eventid="1820" heatid="9430" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:22.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.20" entrycourse="SCM" eventid="1848" heatid="9466" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:22.20" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.16" entrycourse="LCM" eventid="1971" heatid="9488" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:58.16" />
                </ENTRY>
                <ENTRY entrytime="00:04:29.25" entrycourse="LCM" eventid="2103" heatid="9610" lane="3">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-11" name="Erlanger Sparkassen-Cup" qualificationtime="00:04:29.25" />
                </ENTRY>
                <ENTRY entrytime="00:08:58.51" entrycourse="LCM" eventid="2168" heatid="9617" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:08:58.51" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:38.48" eventid="5316" heatid="9481" lane="3">
                  <MEETINFO city="Dachau" date="2019-02-16" name="20. Int. Dachauer Masters-Cup" qualificationtime="00:02:01.52" />
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6143" number="1" />
                    <RELAYPOSITION athleteid="6101" number="2" />
                    <RELAYPOSITION athleteid="6123" number="3" />
                    <RELAYPOSITION athleteid="6097" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY entrytime="00:01:42.14" eventid="2232" heatid="9620" lane="1">
                  <MEETINFO city="Dachau" date="2019-02-17" name="20. Int. Dachauer Masters-Cup" qualificationtime="00:01:54.08" />
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6097" number="1" />
                    <RELAYPOSITION athleteid="6123" number="2" />
                    <RELAYPOSITION athleteid="6155" number="3" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:36.15" eventid="1855" heatid="9477" lane="3">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:42.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.03" eventid="5303" heatid="9615" lane="4">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:55.28" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4328" nation="GER" region="02" clubid="6408" name="SSG Bad Reichenhall im BGL e.V.">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Stephanie" gender="F" lastname="Schneider" nation="GER" license="277641" athleteid="6409">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.25" entrycourse="SCM" eventid="1785" heatid="9399" lane="1">
                  <MEETINFO city="Rosenheim" course="SCM" date="2019-02-09" name="Obb Kreis- und Keisjahrgangsmeisterschaften K 2" qualificationtime="00:01:12.25" />
                </ENTRY>
                <ENTRY entrytime="00:04:55.50" entrycourse="SCM" eventid="5320" heatid="9472" lane="3">
                  <MEETINFO city="Rif" course="SCM" date="2019-02-03" name="Int. Salzburger Kurzbahn Landesmeisterschaft" qualificationtime="00:04:55.50" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.13" entrycourse="SCM" eventid="1978" heatid="9501" lane="1">
                  <MEETINFO city="Rif" course="SCM" date="2019-02-02" name="Int. Salzburger Kurzbahn Landesmeisterschaft" qualificationtime="00:02:20.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.84" entrycourse="SCM" eventid="2075" heatid="9562" lane="2">
                  <MEETINFO city="Rosenheim" course="SCM" date="2019-02-09" name="Obb Kreis- und Keisjahrgangsmeisterschaften K 2" qualificationtime="00:02:38.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6695" nation="GER" region="02" clubid="6942" name="SSG Coburg">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Miklos" gender="M" lastname="Kalocsai" nation="GER" license="350497" athleteid="6943">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.50" entrycourse="SCM" eventid="1778" heatid="9390" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:02.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.19" entrycourse="SCM" eventid="1834" heatid="9447" lane="1">
                  <MEETINFO city="Coburg" course="SCM" date="2019-06-30" name="Stadtmeisterschaft Coburg" qualificationtime="00:00:26.27" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.80" entrycourse="SCM" eventid="2027" heatid="9544" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:05.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.83" entrycourse="SCM" eventid="5307" heatid="9594" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:27.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Hannah" gender="F" lastname="Liebkopf" nation="GER" license="316810" athleteid="6948">
              <ENTRIES>
                <ENTRY entrytime="00:02:33.00" entrycourse="SCM" eventid="1813" heatid="9425" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:30.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.60" entrycourse="SCM" eventid="1841" heatid="9460" lane="4">
                  <MEETINFO city="Coburg" course="LCM" date="2019-05-25" name="41. Jahrgangs- und Pokalschwimmen am 25.05." qualificationtime="00:00:31.25" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.57" entrycourse="SCM" eventid="2006" heatid="9530" lane="1">
                  <MEETINFO city="Coburg" course="SCM" date="2019-06-30" name="Stadtmeisterschaft Coburg" qualificationtime="00:01:07.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.48" entrycourse="SCM" eventid="2075" heatid="9564" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:32.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Carlota" gender="F" lastname="Schmidt-Bäumler Fernández" nation="GER" license="346096" athleteid="6953">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.69" entrycourse="SCM" eventid="1841" heatid="9459" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:30.69" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.73" entrycourse="SCM" eventid="2006" heatid="9528" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:09.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Mia" gender="F" lastname="Teodorovic" nation="GER" license="380176" athleteid="6956">
              <ENTRIES>
                <ENTRY entrytime="00:22:34.17" entrycourse="LCM" eventid="5318" heatid="9478" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-01-19" name="Bayerische Meisterschaften lange Strecken" qualificationtime="00:22:34.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4330" nation="GER" region="02" clubid="6654" name="SSG Neptun Germering">
          <ATHLETES>
            <ATHLETE birthdate="2006-01-01" firstname="Maia" gender="F" lastname="David" nation="GER" license="428978" athleteid="6655">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.36" entrycourse="SCM" eventid="1756" heatid="9371" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:36.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.14" entrycourse="SCM" eventid="2089" heatid="9581" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:29.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Claudia" gender="F" lastname="Dobmeier" nation="GER" license="299888" athleteid="6658">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.36" entrycourse="SCM" eventid="1059" heatid="9346" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:04.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.87" entrycourse="SCM" eventid="2089" heatid="9582" lane="3">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:28.86" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Florian" gender="M" lastname="Dobmeier" nation="GER" license="331618" athleteid="6661">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.43" entrycourse="SCM" eventid="1834" heatid="9445" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:26.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.42" entrycourse="SCM" eventid="1971" heatid="9487" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:58.42" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Niklas" gender="M" lastname="Fink" nation="GER" license="376169" athleteid="6664">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.13" entrycourse="SCM" eventid="1778" heatid="9389" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:03.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.43" entrycourse="SCM" eventid="1834" heatid="9446" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:26.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.84" entrycourse="SCM" eventid="1971" heatid="9486" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:58.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.71" entrycourse="SCM" eventid="5307" heatid="9594" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:27.71" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Florian" gender="M" lastname="Golda" nation="GER" license="371166" athleteid="6669">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.74" entrycourse="SCM" eventid="1985" heatid="9510" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:33.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Johannes" gender="M" lastname="Mais" nation="GER" license="283682" athleteid="6671">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.49" entrycourse="SCM" eventid="1778" heatid="9390" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:02.49" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.83" entrycourse="SCM" eventid="1971" heatid="9488" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:57.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.08" entrycourse="SCM" eventid="5307" heatid="9594" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:28.08" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Lukas" gender="M" lastname="Mais" nation="GER" license="283683" athleteid="6675">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.81" entrycourse="SCM" eventid="1834" heatid="9444" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:26.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.53" entrycourse="SCM" eventid="1971" heatid="9486" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:58.53" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Luis" gender="M" lastname="Obermayer" nation="GER" license="301457" athleteid="6678">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.88" entrycourse="SCM" eventid="1763" heatid="9380" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:10.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.10" entrycourse="SCM" eventid="1820" heatid="9429" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:25.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.18" entrycourse="SCM" eventid="1834" heatid="9442" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:27.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.39" entrycourse="SCM" eventid="1985" heatid="9512" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:32.39" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.65" entrycourse="SCM" eventid="2027" heatid="9542" lane="4">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:01:06.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.15" entrycourse="SCM" eventid="2082" heatid="9572" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:36.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Johannes" gender="M" lastname="Sedlmayer" nation="GER" license="334946" athleteid="6685">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.69" entrycourse="SCM" eventid="1763" heatid="9377" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:14.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.23" entrycourse="SCM" eventid="1985" heatid="9509" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:34.23" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Alessia" gender="F" lastname="Tammaro" nation="GER" license="333921" athleteid="6688">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.87" entrycourse="SCM" eventid="1785" heatid="9398" lane="6">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:01:12.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.36" entrycourse="SCM" eventid="2034" heatid="9551" lane="5">
                  <MEETINFO city="Dachau" course="SCM" date="2019-02-10" name="Kreisjahrgangsmeisterschaften Kreis4 Obb." qualificationtime="00:00:33.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Benedikt" gender="M" lastname="Waechter" nation="GER" license="325820" athleteid="6691">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.18" entrycourse="SCM" eventid="1834" heatid="9442" lane="3">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:27.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.38" entrycourse="SCM" eventid="1971" heatid="9485" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:59.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.00" eventid="1855" heatid="9476" lane="5">
                  <MEETINFO city="Kaufering" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:22.48" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.00" eventid="5303" heatid="9614" lane="6">
                  <MEETINFO city="Pappenheim" date="2019-07-13" name="Bay. Meisterschaften  Masters" qualificationtime="00:02:10.11" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4331" nation="GER" region="02" clubid="5951" name="SSKC Poseidon Aschaffenburg">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Cäcilia" gender="F" lastname="Bausback" nation="GER" license="308503" athleteid="5952">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.37" entrycourse="LCM" eventid="1059" heatid="9350" lane="1">
                  <MEETINFO city="Gzira" course="LCM" date="2019-04-25" name="Easter International Meet" qualificationtime="00:01:03.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.58" entrycourse="SCM" eventid="1813" heatid="9426" lane="2">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-04" name="69.Süddeutsche Meisterschaften" qualificationtime="00:02:27.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.85" entrycourse="LCM" eventid="1841" heatid="9463" lane="5">
                  <MEETINFO city="Gzira" course="LCM" date="2019-04-26" name="Easter International Meet" qualificationtime="00:00:29.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.78" entrycourse="SCM" eventid="2006" heatid="9529" lane="2">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-05" name="69.Süddeutsche Meisterschaften" qualificationtime="00:01:06.78" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.38" entrycourse="SCM" eventid="2096" heatid="9605" lane="1">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:02:31.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Lea" gender="F" lastname="Becker" nation="GER" license="343847" athleteid="5958">
              <ENTRIES>
                <ENTRY entrytime="00:05:37.88" entrycourse="SCM" eventid="1771" heatid="9387" lane="5">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:05:37.88" />
                </ENTRY>
                <ENTRY entrytime="00:04:57.00" entrycourse="SCM" eventid="5320" heatid="9472" lane="5">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-05-31" name="Main-Echo Cup" qualificationtime="00:05:08.17" />
                </ENTRY>
                <ENTRY entrytime="00:20:36.74" entrycourse="SCM" eventid="5318" heatid="9478" lane="4">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:20:36.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.09" entrycourse="SCM" eventid="2034" heatid="9549" lane="3">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:00:34.09" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.31" entrycourse="SCM" eventid="2096" heatid="9603" lane="2">
                  <MEETINFO city="Hofheim am Taunus" course="SCM" date="2019-05-26" name="12. Hofheimer Frühjahrsmeeting" qualificationtime="00:02:35.31" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Carlotta" gender="F" lastname="Fröhlich" nation="GER" license="326201" athleteid="5964">
              <ENTRIES>
                <ENTRY entrytime="00:05:29.40" entrycourse="SCM" eventid="1771" heatid="9388" lane="6">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:05:29.40" />
                </ENTRY>
                <ENTRY entrytime="00:04:57.00" entrycourse="SCM" eventid="5320" heatid="9472" lane="2">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-05-31" name="Main-Echo Cup" qualificationtime="00:05:02.34" />
                </ENTRY>
                <ENTRY entrytime="00:19:53.83" entrycourse="SCM" eventid="5318" heatid="9479" lane="1">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:19:53.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.88" entrycourse="SCM" eventid="1978" heatid="9500" lane="2">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:02:20.88" />
                </ENTRY>
                <ENTRY entrytime="00:10:26.31" entrycourse="SCM" eventid="2020" heatid="9541" lane="1">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:10:26.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.04" entrycourse="SCM" eventid="2089" heatid="9577" lane="1">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:00:30.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Alexander" gender="M" lastname="Gening" nation="GER" license="376694" athleteid="5971">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.58" entrycourse="SCM" eventid="1763" heatid="9377" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:14.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.42" entrycourse="LCM" eventid="1820" heatid="9430" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:23.42" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.66" entrycourse="SCM" eventid="1985" heatid="9510" lane="5">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:00:33.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:39.98" entrycourse="SCM" eventid="2082" heatid="9570" lane="5">
                  <MEETINFO city="Gzira" course="LCM" date="2019-04-26" name="Easter International Meet" qualificationtime="00:02:39.98" />
                </ENTRY>
                <ENTRY entrytime="00:04:35.05" entrycourse="LCM" eventid="2103" heatid="9609" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:35.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1995-01-01" firstname="Nils" gender="M" lastname="Haack" nation="GER" license="265043" athleteid="5977">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.05" entrycourse="LCM" eventid="1749" heatid="9364" lane="5">
                  <MEETINFO city="Gzira" course="LCM" date="2019-04-26" name="Easter International Meet" qualificationtime="00:02:08.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.95" entrycourse="SCM" eventid="1834" heatid="9448" lane="2">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:00:25.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.70" entrycourse="SCM" eventid="1971" heatid="9492" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:55.79" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.56" entrycourse="SCM" eventid="2041" heatid="9559" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:15.19" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Alexander" gender="M" lastname="Hebeler" nation="GER" license="297466" athleteid="5982">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.59" entrycourse="SCM" eventid="1763" heatid="9378" lane="3">
                  <MEETINFO city="Hofheim am Taunus" course="SCM" date="2019-05-26" name="12. Hofheimer Frühjahrsmeeting" qualificationtime="00:01:12.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.66" entrycourse="SCM" eventid="1834" heatid="9444" lane="3">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:00:26.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.89" entrycourse="SCM" eventid="1971" heatid="9486" lane="6">
                  <MEETINFO city="Hofheim am Taunus" course="SCM" date="2019-05-26" name="12. Hofheimer Frühjahrsmeeting" qualificationtime="00:00:58.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.14" entrycourse="SCM" eventid="1985" heatid="9513" lane="1">
                  <MEETINFO city="Hofheim am Taunus" course="SCM" date="2019-05-26" name="12. Hofheimer Frühjahrsmeeting" qualificationtime="00:00:32.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Anika" gender="F" lastname="Heinz" nation="GER" license="316543" athleteid="5987">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.92" entrycourse="SCM" eventid="1059" heatid="9352" lane="3">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:01:00.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.66" entrycourse="SCM" eventid="1785" heatid="9400" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-06" name="Ufr. Langbahn- und 2. int. Mastersmeisterschaften" qualificationtime="00:01:13.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.91" entrycourse="SCM" eventid="1841" heatid="9459" lane="6">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:00:30.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.38" entrycourse="SCM" eventid="2006" heatid="9528" lane="3">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:01:09.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.14" entrycourse="SCM" eventid="2034" heatid="9554" lane="1">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-04-11" name="Landesfinale bay. Schulen JtfO" qualificationtime="00:00:32.14" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.20" entrycourse="SCM" eventid="2089" heatid="9584" lane="4">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-04-11" name="Landesfinale bay. Schulen JtfO" qualificationtime="00:00:28.27" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Fabienne" gender="F" lastname="Krüger" nation="GER" license="297473" athleteid="5994">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.57" entrycourse="SCM" eventid="1059" heatid="9354" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:00.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.35" eventid="1799" heatid="9414" lane="5" />
                <ENTRY entrytime="00:00:30.25" entrycourse="LCM" eventid="1841" heatid="9461" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:31.32" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.25" entrycourse="LCM" eventid="1978" heatid="9505" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:14.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.64" entrycourse="SCM" eventid="2089" heatid="9586" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:27.64" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Hannah" gender="F" lastname="Ludwig" nation="GER" license="314591" athleteid="6000">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.54" entrycourse="SCM" eventid="1756" heatid="9370" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:36.54" />
                </ENTRY>
                <ENTRY entrytime="00:02:54.50" entrycourse="SCM" eventid="1827" heatid="9436" lane="3">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:02:54.50" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.99" entrycourse="SCM" eventid="1992" heatid="9519" lane="4">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:01:20.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.10" entrycourse="SCM" eventid="2089" heatid="9576" lane="4">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:00:30.39" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Anna" gender="F" lastname="Reibenspiess" nation="GER" license="297472" athleteid="6005">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.95" entrycourse="LCM" eventid="1059" heatid="9354" lane="2">
                  <MEETINFO city="Seraing" course="LCM" date="2019-01-27" name="Meeting de Janus" qualificationtime="00:01:00.98" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.09" entrycourse="SCM" eventid="1813" heatid="9426" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:23.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.31" entrycourse="LCM" eventid="1841" heatid="9463" lane="4">
                  <MEETINFO city="Heidelberg" course="LCM" date="2019-03-24" name="Nikar - Cup" qualificationtime="00:00:29.31" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.22" entrycourse="LCM" eventid="2006" heatid="9529" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:01:03.22" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.61" entrycourse="LCM" eventid="2075" heatid="9566" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:22.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Mia-Sophie" gender="F" lastname="Sauer" nation="GER" license="363437" athleteid="6011">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.66" entrycourse="SCM" eventid="1785" heatid="9399" lane="4">
                  <MEETINFO city="Hofheim am Taunus" course="SCM" date="2019-05-26" name="12. Hofheimer Frühjahrsmeeting" qualificationtime="00:01:11.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.00" entrycourse="SCM" eventid="1841" heatid="9457" lane="1">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:00:32.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.08" entrycourse="SCM" eventid="2034" heatid="9551" lane="4">
                  <MEETINFO city="Hofheim am Taunus" course="SCM" date="2019-05-26" name="12. Hofheimer Frühjahrsmeeting" qualificationtime="00:00:33.08" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.15" entrycourse="SCM" eventid="2096" heatid="9606" lane="6">
                  <MEETINFO city="Hofheim am Taunus" course="SCM" date="2019-05-26" name="12. Hofheimer Frühjahrsmeeting" qualificationtime="00:02:33.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Franka" gender="F" lastname="Timm" nation="GER" license="343859" athleteid="6016">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.55" entrycourse="SCM" eventid="1756" heatid="9370" lane="1">
                  <MEETINFO city="Gzira" course="LCM" date="2019-04-25" name="Easter International Meet" qualificationtime="00:00:36.55" />
                </ENTRY>
                <ENTRY entrytime="00:02:55.27" entrycourse="SCM" eventid="1827" heatid="9436" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:55.27" />
                </ENTRY>
                <ENTRY entrytime="00:19:58.95" entrycourse="SCM" eventid="5318" heatid="9479" lane="6">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:19:58.95" />
                </ENTRY>
                <ENTRY entrytime="00:01:19.30" entrycourse="SCM" eventid="1992" heatid="9521" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:19.30" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.21" entrycourse="LCM" eventid="2089" heatid="9580" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:29.21" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2000-01-01" firstname="Philipp" gender="M" lastname="Walter" nation="GER" license="284784" athleteid="6022">
              <ENTRIES>
                <ENTRY entrytime="00:02:17.16" entrycourse="SCM" eventid="1820" heatid="9433" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:17.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.86" entrycourse="SCM" eventid="1848" heatid="9468" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:17.12" />
                </ENTRY>
                <ENTRY entrytime="00:04:54.59" entrycourse="SCM" eventid="1999" heatid="9527" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:04:54.59" />
                </ENTRY>
                <ENTRY entrytime="00:04:23.56" entrycourse="SCM" eventid="2103" heatid="9612" lane="1">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-05-31" name="Main-Echo Cup" qualificationtime="00:04:23.56" />
                </ENTRY>
                <ENTRY entrytime="00:09:06.64" entrycourse="SCM" eventid="2168" heatid="9617" lane="6">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:09:19.45" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Jule" gender="F" lastname="Weindel" nation="GER" license="314609" athleteid="6028">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.77" entrycourse="SCM" eventid="1059" heatid="9351" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:02.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.30" eventid="1799" heatid="9413" lane="6" />
                <ENTRY entrytime="00:00:30.75" entrycourse="LCM" eventid="1841" heatid="9459" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:30.75" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.99" entrycourse="SCM" eventid="1992" heatid="9519" lane="3">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:01:20.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.22" entrycourse="SCM" eventid="2089" heatid="9584" lane="2">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-06-01" name="Main-Echo Cup" qualificationtime="00:00:28.57" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.06" eventid="5314" heatid="9482" lane="4">
                  <MEETINFO city="Gau-Algesheim" date="2019-01-20" name="30. Internationale Masters mit RLP-KBM" qualificationtime="00:02:16.42" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.06" eventid="2224" heatid="9618" lane="5">
                  <MEETINFO city="Gau-Algesheim" date="2019-01-20" name="30. Internationale Masters mit RLP-KBM" qualificationtime="00:02:02.89" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.51" eventid="5303" heatid="9614" lane="1">
                  <MEETINFO city="Gau-Algesheim" date="2019-01-20" name="30. Internationale Masters mit RLP-KBM" qualificationtime="00:02:21.87" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4332" nation="GER" region="02" clubid="6414" name="SSV Forchheim">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Nina" gender="F" lastname="Hohenberger" nation="GER" license="348318" athleteid="6415">
              <ENTRIES>
                <ENTRY entrytime="00:02:36.87" entrycourse="SCM" eventid="2096" heatid="9602" lane="2">
                  <MEETINFO city="Nürnberg" course="LCM" date="2019-07-06" name="Mittelfränkische Meisterschaften" qualificationtime="00:02:41.06" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Lukas" gender="M" lastname="Mursak" nation="GER" license="348315" athleteid="6417">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.63" entrycourse="SCM" eventid="1778" heatid="9390" lane="4">
                  <MEETINFO city="Nürnberg" course="LCM" date="2019-07-06" name="Mittelfränkische Meisterschaften" qualificationtime="00:01:03.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.50" entrycourse="LCM" eventid="1971" heatid="9484" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:00.45" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.30" entrycourse="SCM" eventid="2041" heatid="9558" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:27.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.79" entrycourse="SCM" eventid="5307" heatid="9592" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:28.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Niklas" gender="M" lastname="Schmidt" nation="GER" license="365981" athleteid="6422">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.64" entrycourse="SCM" eventid="1806" heatid="9418" lane="3">
                  <MEETINFO city="Forchheim" course="SCM" date="2019-03-23" name="16. Frühjahrs-Sprint-Meeting_Ausschreibung" qualificationtime="00:00:31.34" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.48" entrycourse="SCM" eventid="1848" heatid="9467" lane="6">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-02-10" name="DMS - , Bezirksliga Mittelfranken" qualificationtime="00:02:21.48" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.39" entrycourse="SCM" eventid="2013" heatid="9534" lane="3">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-02-10" name="DMS - , Bezirksliga Mittelfranken" qualificationtime="00:01:06.79" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4344" nation="GER" region="02" clubid="5739" name="SV Augsburg 1911">
          <ATHLETES>
            <ATHLETE birthdate="1989-01-01" firstname="Nadine" gender="F" lastname="Bender" nation="GER" license="197915" athleteid="5740">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.40" entrycourse="SCM" eventid="1059" heatid="9354" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:00.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.50" entrycourse="SCM" eventid="1785" heatid="9402" lane="1">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:09.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.00" entrycourse="SCM" eventid="1978" heatid="9504" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:13.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.40" eventid="2034" heatid="9553" lane="4" />
                <ENTRY entrytime="00:00:26.97" entrycourse="LCM" eventid="2089" heatid="9586" lane="4">
                  <MEETINFO city="Kempten" course="LCM" date="2019-07-06" name="Bezirksmeisterschaften und Masters" qualificationtime="00:00:29.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1992-01-01" firstname="Matthias" gender="M" lastname="Kopfmüller" nation="GER" license="137031" athleteid="5746">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.61" entrycourse="SCM" eventid="1806" heatid="9420" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:00:28.61" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.90" entrycourse="SCM" eventid="1834" heatid="9453" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:23.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.40" entrycourse="SCM" eventid="1971" heatid="9497" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:00:54.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.40" entrycourse="SCM" eventid="5307" heatid="9594" lane="3">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:27.54" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1977-01-01" firstname="Andreas" gender="M" lastname="Kornes" nation="GER" license="75398" athleteid="5750">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.90" entrycourse="SCM" eventid="1763" heatid="9384" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:05.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.40" entrycourse="SCM" eventid="1834" heatid="9454" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:24.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.50" entrycourse="SCM" eventid="1985" heatid="9516" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:00:29.89" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.00" entrycourse="SCM" eventid="2082" heatid="9573" lane="4">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:24.29" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Robin" gender="M" lastname="Lienhart" nation="GER" license="349208" athleteid="5755">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.62" entrycourse="SCM" eventid="1749" heatid="9361" lane="5">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:05.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.79" entrycourse="SCM" eventid="1834" heatid="9444" lane="1">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:26.79" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.71" entrycourse="SCM" eventid="1848" heatid="9466" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:22.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.18" entrycourse="SCM" eventid="1971" heatid="9487" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:00:58.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.57" entrycourse="SCM" eventid="1985" heatid="9510" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:33.57" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.16" entrycourse="SCM" eventid="2082" heatid="9571" lane="6">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:36.16" />
                </ENTRY>
                <ENTRY entrytime="00:04:25.56" entrycourse="SCM" eventid="2103" heatid="9611" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:04:25.56" />
                </ENTRY>
                <ENTRY entrytime="00:09:10.43" entrycourse="LCM" eventid="2168" heatid="9616" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:09:10.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1989-01-01" firstname="Kornelia" gender="F" lastname="Saal" nation="GER" license="106363" athleteid="5764">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.90" eventid="1756" heatid="9374" lane="5" />
                <ENTRY entrytime="00:01:08.00" eventid="1799" heatid="9413" lane="3" />
                <ENTRY entrytime="00:00:29.50" entrycourse="SCM" eventid="1841" heatid="9461" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:00:29.67" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.50" entrycourse="SCM" eventid="2006" heatid="9529" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:06.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.00" eventid="2075" heatid="9567" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sarah" gender="F" lastname="Sauer" nation="GER" license="342521" athleteid="5770">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.81" entrycourse="SCM" eventid="1059" heatid="9351" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:01.81" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.14" entrycourse="SCM" eventid="1785" heatid="9400" lane="4">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:10.14" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.54" entrycourse="SCM" eventid="1813" heatid="9426" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:27.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.88" entrycourse="SCM" eventid="1841" heatid="9459" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:30.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.78" entrycourse="SCM" eventid="1978" heatid="9503" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:15.78" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.24" entrycourse="SCM" eventid="2006" heatid="9529" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:07.24" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.13" entrycourse="SCM" eventid="2096" heatid="9604" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:29.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1986-01-01" firstname="Matthias" gender="M" lastname="Schwab" nation="GER" license="132395" athleteid="5778">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.90" entrycourse="SCM" eventid="1763" heatid="9382" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:06.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.00" entrycourse="SCM" eventid="1778" heatid="9391" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:59.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.40" entrycourse="SCM" eventid="1985" heatid="9515" lane="4">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:31.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.50" entrycourse="SCM" eventid="5307" heatid="9599" lane="1">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:27.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lux-Sophie" gender="F" lastname="Staudinger" nation="GER" license="354789" athleteid="5783">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.63" entrycourse="SCM" eventid="1059" heatid="9352" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:01.63" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.09" entrycourse="SCM" eventid="1799" heatid="9409" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:13.09" />
                </ENTRY>
                <ENTRY entrytime="00:04:43.26" entrycourse="SCM" eventid="5320" heatid="9474" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:04:43.26" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.25" entrycourse="SCM" eventid="1978" heatid="9504" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:13.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.17" entrycourse="SCM" eventid="2089" heatid="9581" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:29.17" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.98" entrycourse="SCM" eventid="2096" heatid="9602" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:35.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Nele" gender="F" lastname="Stürmer" nation="GER" license="346436" athleteid="5790">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.44" entrycourse="SCM" eventid="1756" heatid="9374" lane="6">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:35.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.79" entrycourse="SCM" eventid="1799" heatid="9408" lane="2">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:14.79" />
                </ENTRY>
                <ENTRY entrytime="00:02:51.72" entrycourse="SCM" eventid="1827" heatid="9437" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:51.72" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.20" entrycourse="SCM" eventid="1992" heatid="9523" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:17.20" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Mark" gender="M" lastname="Toprak" nation="GER" license="346434" athleteid="5795">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.93" entrycourse="SCM" eventid="1763" heatid="9382" lane="4">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:07.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.26" entrycourse="SCM" eventid="1778" heatid="9394" lane="2">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:00:59.18" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.75" entrycourse="SCM" eventid="1834" heatid="9451" lane="3">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:24.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.00" eventid="5316" heatid="9481" lane="2">
                  <MEETINFO city="Augsburg" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:52.44" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.00" eventid="5314" heatid="9483" lane="6">
                  <MEETINFO city="Augsburg" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:06.97" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:43.00" eventid="1855" heatid="9477" lane="2">
                  <MEETINFO city="Augsburg" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:46.23" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.50" eventid="5303" heatid="9615" lane="5">
                  <MEETINFO city="Augsburg" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:56.55" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4347" nation="GER" region="02" clubid="7097" name="SV Bayreuth">
          <ATHLETES>
            <ATHLETE birthdate="1997-01-01" firstname="Sebastian" gender="M" lastname="Feser" nation="GER" license="173941" athleteid="7098">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.12" entrycourse="SCM" eventid="1749" heatid="9363" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:54.93" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.59" entrycourse="SCM" eventid="1778" heatid="9394" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:00:59.94" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.23" entrycourse="SCM" eventid="1820" heatid="9432" lane="4">
                  <MEETINFO city="Pegnitz" course="SCM" date="2019-10-05" name="2. CabrioSol Cup" qualificationtime="00:02:16.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.54" entrycourse="SCM" eventid="1971" heatid="9494" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:53.08" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.01" entrycourse="LCM" eventid="2013" heatid="9536" lane="2">
                  <MEETINFO city="Karlsruhe" course="LCM" date="2019-06-01" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:01:04.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.27" entrycourse="SCM" eventid="5307" heatid="9595" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:00:26.92" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Nico" gender="M" lastname="Heilmann" nation="GER" license="291040" athleteid="7105">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.35" entrycourse="SCM" eventid="1749" heatid="9361" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:02:05.35" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.35" entrycourse="SCM" eventid="1763" heatid="9380" lane="4">
                  <MEETINFO city="Pegnitz" course="SCM" date="2019-10-05" name="2. CabrioSol Cup" qualificationtime="00:01:10.35" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.65" entrycourse="SCM" eventid="1820" heatid="9432" lane="6">
                  <MEETINFO city="Pegnitz" course="SCM" date="2019-10-05" name="2. CabrioSol Cup" qualificationtime="00:02:20.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.25" entrycourse="SCM" eventid="1834" heatid="9447" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:26.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.53" entrycourse="SCM" eventid="1971" heatid="9489" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:57.53" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.21" entrycourse="SCM" eventid="2027" heatid="9543" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:05.21" />
                </ENTRY>
                <ENTRY entrytime="00:04:29.17" entrycourse="SCM" eventid="2103" heatid="9611" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:04:29.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4385" nation="GER" region="02" clubid="7299" name="SV Fürstenfeldbrucker Wasserratten e.V.">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Lara" gender="F" lastname="Fink" nation="GER" license="388898" athleteid="7300">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.99" entrycourse="SCM" eventid="1059" heatid="9346" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:05.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.92" entrycourse="SCM" eventid="2089" heatid="9578" lane="1">
                  <MEETINFO city="Erlangen" course="LCM" date="2019-05-11" name="Erlanger Sparkassen-Cup" qualificationtime="00:00:29.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Miriam" gender="F" lastname="Karcher" nation="GER" license="316822" athleteid="7303">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.35" entrycourse="SCM" eventid="1059" heatid="9348" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:03.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.34" entrycourse="SCM" eventid="1756" heatid="9371" lane="1">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:00:35.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.60" entrycourse="SCM" eventid="1799" heatid="9411" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:11.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.69" entrycourse="SCM" eventid="1841" heatid="9457" lane="4">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:31.22" />
                </ENTRY>
                <ENTRY entrytime="00:01:20.51" entrycourse="SCM" eventid="1992" heatid="9520" lane="5">
                  <MEETINFO city="Dachau" course="SCM" date="2019-02-10" name="Kreisjahrgangsmeisterschaften Kreis4 Obb." qualificationtime="00:01:19.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.72" entrycourse="SCM" eventid="2034" heatid="9550" lane="4">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:33.04" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.78" entrycourse="SCM" eventid="2075" heatid="9563" lane="1">
                  <MEETINFO city="Bad Tölz" course="SCM" date="2019-02-24" name="DMS Bezirksdurchgang Oberbayern" qualificationtime="00:02:38.08" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.01" entrycourse="SCM" eventid="2089" heatid="9581" lane="3">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:28.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Felix" gender="M" lastname="Mende" nation="GER" license="312415" athleteid="7312">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.55" entrycourse="SCM" eventid="1763" heatid="9380" lane="5">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:01:10.80" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.99" entrycourse="SCM" eventid="1834" heatid="9448" lane="5">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:25.99" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Lea" gender="F" lastname="Obermair" nation="GER" license="230355" athleteid="7315">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.11" entrycourse="SCM" eventid="1059" heatid="9350" lane="5">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:01:02.11" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.04" entrycourse="SCM" eventid="1785" heatid="9400" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:10.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Janina" gender="F" lastname="Ruoff" nation="GER" license="345905" athleteid="7318">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.13" entrycourse="SCM" eventid="2034" heatid="9549" lane="4">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:34.13" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Julia" gender="F" lastname="Schober" nation="GER" license="362533" athleteid="7320">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.58" entrycourse="SCM" eventid="1756" heatid="9368" lane="4">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:37.58" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.02" entrycourse="SCM" eventid="2089" heatid="9577" lane="2">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:30.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Corinna" gender="F" lastname="Wirkner" nation="GER" license="344665" athleteid="7323">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.00" entrycourse="SCM" eventid="1059" heatid="9352" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:01.00" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.48" entrycourse="SCM" eventid="1785" heatid="9400" lane="5">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:01:10.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.33" entrycourse="SCM" eventid="1841" heatid="9463" lane="6">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:00:30.03" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.77" entrycourse="SCM" eventid="1978" heatid="9503" lane="2">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-06" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:02:15.77" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.83" entrycourse="SCM" eventid="2034" heatid="9552" lane="5">
                  <MEETINFO city="Karlsfeld" course="SCM" date="2019-05-18" name="Kreissprint &amp; Lange Kreis 4 Obb" qualificationtime="00:00:32.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.55" entrycourse="SCM" eventid="2089" heatid="9588" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:27.55" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:01:48.00" eventid="2224" heatid="9618" lane="3">
                  <MEETINFO city="Kaufering" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:01:47.80" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.00" eventid="5314" heatid="9483" lane="3" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4356" nation="GER" region="02" clubid="5541" name="SV GR.-W. Holzkirchen">
          <ATHLETES>
            <ATHLETE birthdate="1996-01-01" firstname="Ludwig" gender="M" lastname="Huber" nation="GER" license="181978" athleteid="5542">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.17" entrycourse="SCM" eventid="1749" heatid="9363" lane="5">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-09" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:02:01.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.45" entrycourse="SCM" eventid="1834" heatid="9452" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-02-09" name="Kreiskurzbahnmeisterschaften K3 Obb." qualificationtime="00:00:24.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.81" entrycourse="SCM" eventid="1971" heatid="9495" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-02-09" name="Kreiskurzbahnmeisterschaften K3 Obb." qualificationtime="00:00:53.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.04" entrycourse="SCM" eventid="5307" heatid="9596" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-02-09" name="Kreiskurzbahnmeisterschaften K3 Obb." qualificationtime="00:00:27.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Moritz" gender="M" lastname="Werner" nation="GER" license="292813" athleteid="5547">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.59" entrycourse="SCM" eventid="1763" heatid="9381" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:08.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.47" entrycourse="SCM" eventid="1834" heatid="9449" lane="4">
                  <MEETINFO city="Kaufbeuren" course="SCM" date="2019-03-23" name="18. Internationaler Buron Cup" qualificationtime="00:00:25.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.84" entrycourse="SCM" eventid="1985" heatid="9514" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:30.52" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.27" entrycourse="SCM" eventid="2027" heatid="9546" lane="6">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:04.27" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.09" entrycourse="SCM" eventid="5307" heatid="9596" lane="6">
                  <MEETINFO city="Kaufbeuren" course="SCM" date="2019-03-24" name="18. Internationaler Buron Cup" qualificationtime="00:00:27.09" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4357" nation="GER" region="02" clubid="5698" name="SV Grafing-Ebersberg">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Amelie" gender="F" lastname="Kiermeier" nation="GER" license="346582" athleteid="6037">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.01" entrycourse="SCM" eventid="1059" heatid="9348" lane="5">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:03.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.38" entrycourse="SCM" eventid="1841" heatid="9462" lane="6">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:30.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Florian" gender="M" lastname="Kühn" nation="GER" license="279242" athleteid="6040">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.85" entrycourse="SCM" eventid="1778" heatid="9392" lane="6">
                  <MEETINFO city="Wetzlar" course="LCM" date="2019-05-04" name="27. Süddeutsche Jahrgangsmeisterschaften" qualificationtime="00:00:59.02" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.26" entrycourse="SCM" eventid="1806" heatid="9420" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:29.39" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.28" entrycourse="SCM" eventid="1848" heatid="9469" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:16.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.86" entrycourse="SCM" eventid="2013" heatid="9538" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:03.37" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.22" entrycourse="SCM" eventid="2041" heatid="9558" lane="2">
                  <MEETINFO city="Wetzlar" course="LCM" date="2019-05-05" name="27. Süddeutsche Jahrgangsmeisterschaften" qualificationtime="00:02:12.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.65" entrycourse="SCM" eventid="5307" heatid="9597" lane="1">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:26.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Silvia" gender="F" lastname="Kühn" nation="GER" license="300827" athleteid="6047">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.57" entrycourse="SCM" eventid="1059" heatid="9352" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:01.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.17" entrycourse="SCM" eventid="1785" heatid="9399" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:11.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.20" entrycourse="SCM" eventid="1841" heatid="9463" lane="1">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:30.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.11" entrycourse="SCM" eventid="2006" heatid="9531" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:08.11" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.24" entrycourse="SCM" eventid="2034" heatid="9555" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:32.24" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.32" entrycourse="SCM" eventid="2089" heatid="9584" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:28.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Luisa" gender="F" lastname="Rumler" nation="GER" license="350378" athleteid="5699">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.74" entrycourse="SCM" eventid="1059" heatid="9351" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:01:00.91" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.81" entrycourse="SCM" eventid="1785" heatid="9401" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:09.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.09" entrycourse="SCM" eventid="1841" heatid="9462" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:29.81" />
                </ENTRY>
                <ENTRY entrytime="00:04:41.11" entrycourse="LCM" eventid="5320" heatid="9474" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:42.70" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.59" entrycourse="SCM" eventid="1978" heatid="9504" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:12.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.51" entrycourse="SCM" eventid="2034" heatid="9552" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:32.44" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.72" entrycourse="SCM" eventid="2075" heatid="9566" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:31.72" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.87" entrycourse="SCM" eventid="2089" heatid="9585" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:27.60" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.93" entrycourse="LCM" eventid="2096" heatid="9605" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:33.93" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.00" entrycourse="SCM" eventid="1799" heatid="9415" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:09.00" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5713" nation="GER" region="02" clubid="5880" name="SV Hengersberg">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Lukas" gender="M" lastname="Eisenschink" nation="GER" license="326212" athleteid="5881">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.04" entrycourse="SCM" eventid="1806" heatid="9418" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:31.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.59" entrycourse="SCM" eventid="1834" heatid="9445" lane="1">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:26.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.41" entrycourse="SCM" eventid="1971" heatid="9489" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:57.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.80" entrycourse="SCM" eventid="2027" heatid="9542" lane="2">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:01:06.85" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Barbara" gender="F" lastname="Leitl" nation="GER" license="310921" athleteid="5886">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.46" entrycourse="SCM" eventid="2089" heatid="9579" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:29.46" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Leo" gender="M" lastname="Loibl" nation="GER" license="357942" athleteid="5888">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.88" entrycourse="SCM" eventid="1834" heatid="9443" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:26.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Erik" gender="M" lastname="Stögbauer" nation="GER" license="291450" athleteid="5890">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.25" entrycourse="SCM" eventid="1834" heatid="9450" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:25.74" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4341" nation="GER" region="02" clubid="5828" name="SV Hof 1911 e. V.">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Marlon" gender="M" lastname="Meisel" nation="GER" license="291289" athleteid="5829">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.69" entrycourse="SCM" eventid="1778" heatid="9392" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:59.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.57" entrycourse="SCM" eventid="1806" heatid="9422" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:27.57" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.12" entrycourse="SCM" eventid="1834" heatid="9450" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2019-10-12" name="Oberfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:25.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.33" entrycourse="SCM" eventid="1971" heatid="9493" lane="4">
                  <MEETINFO city="Plauen" course="SCM" date="2019-09-28" name="Plauener Herbst-Mehrkampf" qualificationtime="00:00:55.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.17" entrycourse="SCM" eventid="2013" heatid="9538" lane="5">
                  <MEETINFO city="Plauen" course="SCM" date="2019-09-28" name="Plauener Herbst-Mehrkampf" qualificationtime="00:01:01.17" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.47" entrycourse="SCM" eventid="5307" heatid="9598" lane="4">
                  <MEETINFO city="Plauen" course="SCM" date="2019-09-28" name="Plauener Herbst-Mehrkampf" qualificationtime="00:00:25.47" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4360" nation="GER" region="02" clubid="6486" name="SV Lohhof">
          <ATHLETES>
            <ATHLETE birthdate="1998-01-01" firstname="Caroline" gender="F" lastname="Titze" nation="GER" license="198707" athleteid="6487">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.84" entrycourse="SCM" eventid="1799" heatid="9413" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:08.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.49" entrycourse="SCM" eventid="1841" heatid="9462" lane="4">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-30" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:29.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.07" entrycourse="LCM" eventid="2006" heatid="9529" lane="1">
                  <MEETINFO city="Heidenheim" course="LCM" date="2019-03-23" name="Internationales Schwimmfest Heidenheim" qualificationtime="00:01:08.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.96" entrycourse="SCM" eventid="2034" heatid="9554" lane="5">
                  <MEETINFO city="Landau/Isar" course="SCM" date="2019-06-29" name="21. Internationales Landauer Sprinter-Treffen" qualificationtime="00:00:31.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.75" entrycourse="SCM" eventid="2089" heatid="9587" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:27.75" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4364" nation="GER" region="02" clubid="6205" name="SV Ottobrunn 1970 e.V.">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Leon" gender="M" lastname="Haslinger" nation="GER" license="316236" athleteid="6206">
              <ENTRIES>
                <ENTRY entrytime="00:18:40.73" eventid="1792" heatid="9406" lane="1" />
                <ENTRY entrytime="00:09:45.19" eventid="2168" status="RJC" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lana" gender="F" lastname="Kreppenhofer" nation="GER" license="345306" athleteid="6209">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.66" entrycourse="SCM" eventid="1059" heatid="9346" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:04.66" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.04" entrycourse="SCM" eventid="1785" heatid="9397" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:13.04" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.76" entrycourse="SCM" eventid="1841" heatid="9457" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:31.76" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.52" entrycourse="SCM" eventid="2075" heatid="9562" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:38.52" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.54" entrycourse="SCM" eventid="2096" heatid="9603" lane="5">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:37.52" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Kenneth" gender="M" lastname="Münster" nation="GER" license="349589" athleteid="6215">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.31" entrycourse="SCM" eventid="1749" heatid="9360" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:07.31" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.23" entrycourse="SCM" eventid="1820" heatid="9429" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:02:26.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.97" entrycourse="SCM" eventid="1834" heatid="9443" lane="2">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:26.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.69" entrycourse="SCM" eventid="1971" heatid="9488" lane="3">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:57.69" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Marlene" gender="F" lastname="Ruf" nation="GER" license="345302" athleteid="6220">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.85" entrycourse="SCM" eventid="1756" heatid="9372" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:34.85" />
                </ENTRY>
                <ENTRY entrytime="00:01:11.15" eventid="1799" heatid="9411" lane="2" />
                <ENTRY entrytime="00:02:46.22" entrycourse="SCM" eventid="1827" heatid="9437" lane="4">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:46.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.88" entrycourse="SCM" eventid="1841" heatid="9459" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:30.88" />
                </ENTRY>
                <ENTRY entrytime="00:01:16.26" entrycourse="SCM" eventid="1992" heatid="9524" lane="5">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-05" name="69.Süddeutsche Meisterschaften" qualificationtime="00:01:16.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.53" entrycourse="SCM" eventid="2006" heatid="9528" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:09.53" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.80" entrycourse="SCM" eventid="2075" heatid="9563" lane="3">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:34.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.61" entrycourse="SCM" eventid="2089" heatid="9578" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:29.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Luisa" gender="F" lastname="Schmitz" nation="GER" license="362017" athleteid="6229">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.08" entrycourse="SCM" eventid="1059" heatid="9345" lane="4">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:05.08" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.30" entrycourse="SCM" eventid="1785" heatid="9397" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:13.30" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lorie" gender="F" lastname="Seranski" nation="GER" license="316888" athleteid="6232">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.65" entrycourse="SCM" eventid="1059" heatid="9353" lane="6">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:01:00.65" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.37" entrycourse="SCM" eventid="1785" heatid="9403" lane="2">
                  <MEETINFO city="Freiburg" course="LCM" date="2019-05-05" name="69.Süddeutsche Meisterschaften" qualificationtime="00:01:06.29" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.96" entrycourse="SCM" eventid="1799" heatid="9415" lane="6">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:09.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.23" entrycourse="SCM" eventid="2034" heatid="9554" lane="4">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:31.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.71" entrycourse="SCM" eventid="2089" heatid="9588" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:27.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.76" entrycourse="SCM" eventid="2096" heatid="9606" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:26.76" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Viet Nghia" gender="M" lastname="Truong" nation="GER" license="311579" athleteid="6239">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.47" entrycourse="SCM" eventid="1763" heatid="9379" lane="6">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:12.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.67" entrycourse="SCM" eventid="1834" heatid="9444" lane="4">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:26.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.54" eventid="1855" heatid="9476" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="6215" number="1" />
                    <RELAYPOSITION number="2" />
                    <RELAYPOSITION athleteid="6232" number="3" />
                    <RELAYPOSITION athleteid="6220" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4384" nation="GER" region="02" clubid="7332" name="SV Wacker Burghausen">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Marie-Therese" gender="F" lastname="Bartl" nation="GER" license="296587" athleteid="7333">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.88" entrycourse="SCM" eventid="1059" heatid="9346" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:02.29" />
                </ENTRY>
                <ENTRY entrytime="00:05:30.56" entrycourse="LCM" eventid="1771" heatid="9387" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-15" name="10. Internationales Frühjahresmeeting" qualificationtime="00:05:30.56" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.47" entrycourse="SCM" eventid="1813" heatid="9426" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:33.47" />
                </ENTRY>
                <ENTRY entrytime="00:04:45.84" entrycourse="SCM" eventid="5320" heatid="9474" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:04:40.07" />
                </ENTRY>
                <ENTRY entrytime="00:18:41.33" entrycourse="LCM" eventid="5318" heatid="9479" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-15" name="10. Internationales Frühjahresmeeting" qualificationtime="00:18:41.33" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Nico" gender="M" lastname="Basten" nation="GER" license="321160" athleteid="7339">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.01" entrycourse="SCM" eventid="1749" heatid="9363" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:02.02" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.90" entrycourse="LCM" eventid="1778" heatid="9389" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-16" name="10. Internationales Frühjahresmeeting" qualificationtime="00:01:06.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.87" entrycourse="SCM" eventid="1806" heatid="9419" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:28.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.60" entrycourse="SCM" eventid="1848" heatid="9468" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:11.60" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.61" entrycourse="LCM" eventid="1971" heatid="9493" lane="1">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:55.61" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.01" entrycourse="SCM" eventid="2013" heatid="9536" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:01:02.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.59" entrycourse="SCM" eventid="5307" heatid="9592" lane="4">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:28.59" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Yannick" gender="M" lastname="Buschhardt" nation="GER" license="227101" athleteid="7347">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.74" entrycourse="SCM" eventid="1806" heatid="9422" lane="2">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:27.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.40" entrycourse="SCM" eventid="1848" heatid="9468" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:08.40" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.60" entrycourse="SCM" eventid="1971" heatid="9491" lane="5">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:57.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.02" entrycourse="SCM" eventid="2013" heatid="9536" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:58.93" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Nicole" gender="F" lastname="Fritsch" nation="GER" license="333674" athleteid="7352">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.30" entrycourse="SCM" eventid="1059" heatid="9355" lane="5">
                  <MEETINFO city="Erding" course="LCM" date="2019-07-06" name="Oberbayerische Jahrgangsmeisterschaften" qualificationtime="00:00:59.64" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.10" entrycourse="SCM" eventid="1785" heatid="9401" lane="2">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:01:07.45" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.10" entrycourse="SCM" eventid="1841" heatid="9461" lane="3">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:29.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Maximilian" gender="M" lastname="Kapsegger" nation="GER" license="321145" athleteid="7356">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.66" entrycourse="SCM" eventid="1763" heatid="9377" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:13.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.87" entrycourse="LCM" eventid="1985" heatid="9511" lane="5">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:32.87" />
                </ENTRY>
                <ENTRY entrytime="00:02:41.85" entrycourse="LCM" eventid="2082" heatid="9570" lane="1">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:02:41.85" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Dominik" gender="M" lastname="Kohlschmid" nation="GER" license="242746" athleteid="7360">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.99" entrycourse="LCM" eventid="1763" heatid="9383" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-05-26" name="Deutsche Hochschulmeisterschaften" qualificationtime="00:01:08.99" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.89" entrycourse="SCM" eventid="1834" heatid="9454" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:23.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.89" entrycourse="LCM" eventid="1985" heatid="9516" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-05-24" name="Deutsche Hochschulmeisterschaften" qualificationtime="00:00:30.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.14" entrycourse="LCM" eventid="5307" heatid="9597" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-05-25" name="Deutsche Hochschulmeisterschaften" qualificationtime="00:00:26.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Manuel" gender="M" lastname="Kohlschmid" nation="GER" license="297980" athleteid="7365">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.12" entrycourse="SCM" eventid="1763" heatid="9383" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:04.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.66" entrycourse="SCM" eventid="1834" heatid="9454" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:23.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.39" entrycourse="SCM" eventid="1971" heatid="9497" lane="2">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:52.39" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.75" entrycourse="SCM" eventid="1985" heatid="9515" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:29.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.14" entrycourse="SCM" eventid="2027" heatid="9545" lane="3">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:59.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Verena" gender="F" lastname="Reisegast" nation="GER" license="326167" athleteid="7371">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.63" entrycourse="SCM" eventid="1059" heatid="9351" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:01.24" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.07" entrycourse="SCM" eventid="1799" heatid="9410" lane="4">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:12.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.68" entrycourse="SCM" eventid="1841" heatid="9457" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:31.68" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.48" entrycourse="SCM" eventid="1978" heatid="9505" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:14.48" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.20" entrycourse="SCM" eventid="2034" heatid="9549" lane="2">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:34.20" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.07" entrycourse="SCM" eventid="2089" heatid="9585" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:28.07" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Paulina" gender="F" lastname="Sandner" nation="GER" license="316586" athleteid="7378">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.92" entrycourse="SCM" eventid="1059" heatid="9351" lane="6">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:00.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.77" entrycourse="SCM" eventid="1756" heatid="9373" lane="2">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:34.77" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.00" entrycourse="SCM" eventid="1799" heatid="9415" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:09.33" />
                </ENTRY>
                <ENTRY entrytime="00:01:15.97" entrycourse="SCM" eventid="1992" heatid="9522" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:15.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.47" entrycourse="SCM" eventid="2075" heatid="9566" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:27.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.17" entrycourse="SCM" eventid="2089" heatid="9584" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-05" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:28.17" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Denis" gender="M" lastname="Sczesny" nation="GER" license="350186" athleteid="7385">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.10" entrycourse="SCM" eventid="1763" heatid="9382" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:08.28" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.50" entrycourse="SCM" eventid="1985" heatid="9514" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:30.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:28.10" entrycourse="SCM" eventid="2082" heatid="9571" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:29.03" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Marlene" gender="F" lastname="Sommoggy von" nation="GER" license="304160" athleteid="7389">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.88" entrycourse="LCM" eventid="1756" heatid="9374" lane="4">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:33.88" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.46" entrycourse="SCM" eventid="1827" heatid="9439" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:36.46" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.56" entrycourse="SCM" eventid="1992" heatid="9523" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:12.66" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.87" entrycourse="SCM" eventid="2075" heatid="9567" lane="2">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:26.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.95" entrycourse="SCM" eventid="2089" heatid="9585" lane="2">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:27.95" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.00" eventid="5316" heatid="9481" lane="1" />
                <ENTRY entrytime="00:01:45.00" eventid="2232" heatid="9619" lane="4" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.00" eventid="5314" heatid="9483" lane="1" />
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.00" eventid="1855" heatid="9477" lane="1">
                  <MEETINFO city="Neuötting" date="2019-04-06" name="2. Altöttinger Nachwuchsschwimmen" qualificationtime="00:02:34.28" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.00" eventid="5303" heatid="9615" lane="1">
                  <MEETINFO city="Neuötting" date="2019-04-06" name="2. Altöttinger Nachwuchsschwimmen" qualificationtime="00:02:44.00" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4387" nation="GER" region="02" clubid="5899" name="SV Weiden">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Linus" gender="M" lastname="Brandl" nation="GER" license="317188" athleteid="5900">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.82" entrycourse="SCM" eventid="1806" heatid="9419" lane="5">
                  <MEETINFO city="Berlin" course="SCM" date="2019-09-25" name="Jugend trainiert für Olympia" qualificationtime="00:00:29.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.32" entrycourse="SCM" eventid="1834" heatid="9446" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:26.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.35" entrycourse="SCM" eventid="1971" heatid="9487" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:58.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.76" entrycourse="SCM" eventid="1985" heatid="9511" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:32.76" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Noah" gender="M" lastname="Brandl" nation="GER" license="300722" athleteid="5905">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.73" entrycourse="SCM" eventid="1778" heatid="9393" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:00.73" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.47" entrycourse="SCM" eventid="1806" heatid="9419" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:00:29.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.54" entrycourse="SCM" eventid="1834" heatid="9445" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:26.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.21" entrycourse="SCM" eventid="1971" heatid="9490" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:57.21" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.22" entrycourse="SCM" eventid="5307" heatid="9595" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:27.22" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Leon" gender="M" lastname="Ducheck" nation="GER" license="317126" athleteid="6896">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.22" entrycourse="SCM" eventid="1763" heatid="9378" lane="5">
                  <MEETINFO city="Tirschenreuth" course="SCM" date="2019-04-28" name="17. Internationale Frühlingsschwimmen mit kindgere" qualificationtime="00:01:13.22" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.74" entrycourse="SCM" eventid="1971" heatid="9484" lane="2">
                  <MEETINFO city="Tirschenreuth" course="SCM" date="2019-02-17" name="Bezirk-Mehrkampfmeisterschaften" qualificationtime="00:00:59.74" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.91" entrycourse="SCM" eventid="1985" heatid="9511" lane="1">
                  <MEETINFO city="Tirschenreuth" course="SCM" date="2019-04-28" name="17. Internationale Frühlingsschwimmen mit kindgere" qualificationtime="00:00:32.91" />
                </ENTRY>
                <ENTRY entrytime="00:02:38.93" entrycourse="LCM" eventid="2082" heatid="9570" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:38.93" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Maxine" gender="F" lastname="Edl" nation="GER" license="322620" athleteid="5911">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.36" entrycourse="SCM" eventid="1785" heatid="9397" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:01:13.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.73" entrycourse="SCM" eventid="2034" heatid="9550" lane="2">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:33.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Alexander" gender="M" lastname="Engel" nation="GER" license="336633" athleteid="5914">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.62" eventid="1763" heatid="9378" lane="4" />
                <ENTRY entrytime="00:00:30.23" entrycourse="SCM" eventid="1806" heatid="9419" lane="6">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-03-17" name="10. Internationales Frühjahresmeeting" qualificationtime="00:00:30.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.98" entrycourse="SCM" eventid="1834" heatid="9451" lane="1">
                  <MEETINFO city="Berlin" course="SCM" date="2019-09-24" name="Jugend trainiert für Olympia" qualificationtime="00:00:24.96" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.23" entrycourse="SCM" eventid="1971" heatid="9494" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:54.23" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.11" entrycourse="SCM" eventid="1985" heatid="9513" lane="5">
                  <MEETINFO city="Berlin" course="SCM" date="2019-09-24" name="Jugend trainiert für Olympia" qualificationtime="00:00:31.99" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.02" entrycourse="SCM" eventid="2027" heatid="9546" lane="1">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:01:04.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Jonas" gender="M" lastname="Gießübl" nation="GER" license="331991" athleteid="5921">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.98" entrycourse="SCM" eventid="1834" heatid="9443" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:26.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.19" entrycourse="SCM" eventid="1985" heatid="9509" lane="4">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:34.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.97" entrycourse="SCM" eventid="5307" heatid="9591" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:28.97" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Benjamin" gender="M" lastname="Schindler" nation="GER" license="377803" athleteid="5925">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.03" entrycourse="SCM" eventid="1749" heatid="9359" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-01-12" name="Bezirk-Kurzbahnmeisterschaften" qualificationtime="00:02:09.03" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.42" entrycourse="SCM" eventid="1834" heatid="9446" lane="5">
                  <MEETINFO city="Berlin" course="SCM" date="2019-09-24" name="Jugend trainiert für Olympia" qualificationtime="00:00:25.98" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.10" entrycourse="SCM" eventid="1971" heatid="9490" lane="5">
                  <MEETINFO city="Weiden" course="SCM" date="2019-10-12" name="Oberpfalz-Wintermeisterschaften" qualificationtime="00:00:57.10" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Moritz" gender="M" lastname="Staudinger" nation="GER" license="341208" athleteid="5929">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.12" entrycourse="SCM" eventid="1763" heatid="9382" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:09.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.15" entrycourse="SCM" eventid="1985" heatid="9515" lane="1">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:31.15" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.00" eventid="5316" heatid="9480" lane="2">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:02:02.82" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.00" eventid="2232" heatid="9619" lane="3">
                  <MEETINFO city="Fürth" date="2019-03-16" name="Bay. Kurzbahnmeisterschaften der Masters" qualificationtime="00:01:48.43" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4339" nation="GER" region="02" clubid="7086" name="SV Würzburg 05">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Tabea" gender="F" lastname="Bär" nation="GER" license="302416" athleteid="7087">
              <ENTRIES>
                <ENTRY entrytime="00:02:37.42" entrycourse="SCM" eventid="2075" heatid="9563" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-07" name="Ufr. Langbahn- und 2. int. Mastersmeisterschaften" qualificationtime="00:02:40.36" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.79" entrycourse="SCM" eventid="2089" heatid="9578" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-07" name="Ufr. Langbahn- und 2. int. Mastersmeisterschaften" qualificationtime="00:00:29.66" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Lisa" gender="F" lastname="Gotthardt" nation="GER" license="325565" athleteid="7090">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.43" entrycourse="SCM" eventid="1785" heatid="9399" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:12.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.38" entrycourse="SCM" eventid="1841" heatid="9461" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:30.38" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Olivia" gender="F" lastname="Lang" nation="GER" license="400833" athleteid="7093">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.60" entrycourse="SCM" eventid="1756" heatid="9368" lane="2">
                  <MEETINFO city="Kleinostheim" course="LCM" date="2019-05-05" name="Nationales Schwimm-Meeting" qualificationtime="00:00:37.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:56.18" entrycourse="SCM" eventid="1827" heatid="9436" lane="1">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-07" name="Ufr. Langbahn- und 2. int. Mastersmeisterschaften" qualificationtime="00:02:56.18" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4405" nation="GER" region="02" clubid="5868" name="TSG Kleinostheim">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Joshua" gender="M" lastname="Jankowski" nation="GER" license="309285" athleteid="5869">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.69" entrycourse="SCM" eventid="1985" heatid="9510" lane="1">
                  <MEETINFO city="Esbjerg" course="SCM" date="2019-05-31" name="22th Danish Swim Cup" qualificationtime="00:00:33.69" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Tim" gender="M" lastname="Krenz" nation="GER" license="289249" athleteid="5871">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.56" entrycourse="SCM" eventid="1763" heatid="9380" lane="1">
                  <MEETINFO city="Esbjerg" course="SCM" date="2019-06-02" name="22th Danish Swim Cup" qualificationtime="00:01:10.56" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.13" entrycourse="SCM" eventid="1971" heatid="9488" lane="1">
                  <MEETINFO city="Esbjerg" course="SCM" date="2019-06-02" name="22th Danish Swim Cup" qualificationtime="00:00:58.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.53" entrycourse="SCM" eventid="1985" heatid="9511" lane="3">
                  <MEETINFO city="Esbjerg" course="SCM" date="2019-05-31" name="22th Danish Swim Cup" qualificationtime="00:00:32.53" />
                </ENTRY>
                <ENTRY entrytime="00:02:35.04" entrycourse="SCM" eventid="2082" heatid="9572" lane="1">
                  <MEETINFO city="Esbjerg" course="SCM" date="2019-06-01" name="22th Danish Swim Cup" qualificationtime="00:02:35.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Chantal" gender="F" lastname="Münch" nation="GER" license="374586" athleteid="5876">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.55" entrycourse="SCM" eventid="2034" heatid="9555" lane="2">
                  <MEETINFO city="Aschaffenburg" course="SCM" date="2019-10-12" name="Rhein-Main Mixed-Challenge" qualificationtime="00:00:32.02" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6655" nation="GER" region="02" clubid="5892" name="TSG Nürnberg">
          <ATHLETES>
            <ATHLETE birthdate="2006-01-01" firstname="Lea" gender="F" lastname="Dreykorn" nation="GER" license="331327" athleteid="5893">
              <ENTRIES>
                <ENTRY entrytime="00:02:52.37" entrycourse="SCM" eventid="1827" heatid="9438" lane="6">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:52.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Tim" gender="M" lastname="Fischer" nation="GER" license="402186" athleteid="5895">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.69" entrycourse="SCM" eventid="1834" heatid="9444" lane="2">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:26.69" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.69" entrycourse="SCM" eventid="1971" heatid="9484" lane="4">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:59.54" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Donald" gender="M" lastname="Forster" nation="GER" license="313606" athleteid="5897">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.26" entrycourse="SCM" eventid="1763" heatid="9378" lane="1">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:01:14.44" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.25" entrycourse="SCM" eventid="1985" heatid="9513" lane="6">
                  <MEETINFO city="Erlangen" course="SCM" date="2019-10-13" name="Mittelfränkische Kurzbahnmeisterschaften" qualificationtime="00:00:32.35" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4407" nation="GER" region="02" clubid="5515" name="TSG Stadtbergen 1892">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Katharina" gender="F" lastname="Jawny" nation="GER" license="339031" athleteid="5516">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.76" entrycourse="SCM" eventid="1059" heatid="9347" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:03.76" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.75" entrycourse="SCM" eventid="1799" heatid="9408" lane="4">
                  <MEETINFO city="Stadtbergen" course="SCM" date="2019-04-28" name="Stadtberger Mehrkampftag" qualificationtime="00:01:14.75" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.35" entrycourse="SCM" eventid="2089" heatid="9579" lane="3">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-10" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:00:29.35" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4411" nation="GER" region="02" clubid="5836" name="TSV 1847 Weilheim">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Lukas" gender="M" lastname="Parockinger" nation="GER" license="339098" athleteid="5837">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.25" entrycourse="SCM" eventid="1749" heatid="9360" lane="3">
                  <MEETINFO city="Kaufbeuren" course="SCM" date="2019-03-23" name="18. Internationaler Buron Cup" qualificationtime="00:02:06.25" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.62" entrycourse="SCM" eventid="1778" heatid="9390" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:01:01.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.01" entrycourse="SCM" eventid="1834" heatid="9448" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:26.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.39" entrycourse="SCM" eventid="1971" heatid="9489" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:56.71" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.84" entrycourse="SCM" eventid="2041" heatid="9558" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:20.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.95" entrycourse="SCM" eventid="5307" heatid="9594" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:27.84" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4413" nation="GER" region="02" clubid="5934" name="TSV 1860 Rosenheim">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Sebastian" gender="M" lastname="Hörnig" nation="GER" license="285006" athleteid="5935">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.53" entrycourse="LCM" eventid="1749" heatid="9361" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:05.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.19" entrycourse="SCM" eventid="1806" heatid="9421" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:29.19" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.83" entrycourse="SCM" eventid="1834" heatid="9449" lane="6">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:25.74" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.55" entrycourse="SCM" eventid="1848" heatid="9466" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:21.55" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.26" entrycourse="SCM" eventid="1971" heatid="9492" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:56.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.41" entrycourse="SCM" eventid="2013" heatid="9535" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:03.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.28" entrycourse="SCM" eventid="5307" heatid="9593" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:28.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Maria" gender="F" lastname="Lengauer" nation="GER" license="319637" athleteid="5943">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.48" entrycourse="SCM" eventid="2089" heatid="9579" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:29.48" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Junchi" gender="M" lastname="Weng" nation="GER" license="397184" athleteid="5945">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.64" entrycourse="SCM" eventid="1749" heatid="9361" lane="1">
                  <MEETINFO city="Rosenheim" course="SCM" date="2019-02-09" name="Obb Kreis- und Keisjahrgangsmeisterschaften K 2" qualificationtime="00:02:05.64" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.41" entrycourse="SCM" eventid="1806" heatid="9421" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:29.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.83" entrycourse="SCM" eventid="1834" heatid="9451" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:24.83" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.47" entrycourse="SCM" eventid="1971" heatid="9494" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:54.47" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.70" entrycourse="SCM" eventid="5307" heatid="9599" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:26.70" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4417" nation="GER" region="02" clubid="5529" name="TSV 1862 Friedberg">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Thomas" gender="M" lastname="Schmeikal" nation="GER" license="322956" athleteid="5530">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.29" entrycourse="SCM" eventid="1763" heatid="9379" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:11.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.82" entrycourse="SCM" eventid="1834" heatid="9443" lane="3">
                  <MEETINFO city="Obergünzburg" course="SCM" date="2019-05-04" name="28. Obergünzburger Schwimmfest" qualificationtime="00:00:26.82" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.41" entrycourse="SCM" eventid="1971" heatid="9487" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:00:58.41" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.27" entrycourse="SCM" eventid="1985" heatid="9509" lane="5">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:33.44" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.78" entrycourse="SCM" eventid="2027" heatid="9543" lane="6">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:05.78" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.98" entrycourse="SCM" eventid="5307" heatid="9591" lane="2">
                  <MEETINFO city="Obergünzburg" course="SCM" date="2019-05-04" name="28. Obergünzburger Schwimmfest" qualificationtime="00:00:28.98" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1998-01-01" firstname="Simon" gender="M" lastname="Stengl" nation="GER" license="250031" athleteid="5537">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.37" entrycourse="SCM" eventid="1834" heatid="9450" lane="6">
                  <MEETINFO city="Gersthofen" course="SCM" date="2019-03-10" name="12. Internationaler Cool-Swimming-Cup" qualificationtime="00:00:25.59" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.32" entrycourse="SCM" eventid="1971" heatid="9493" lane="3">
                  <MEETINFO city="Immenstadt" course="SCM" date="2019-02-10" name="DMS, Bezirksliga Schwaben" qualificationtime="00:00:55.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.85" entrycourse="SCM" eventid="2013" heatid="9536" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-03-17" name="Regionalen Bestenkämpfe  - Region Nord" qualificationtime="00:01:02.85" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4445" nation="GER" region="02" clubid="6405" name="TSV 1909 Gersthofen">
          <ATHLETES>
            <ATHLETE birthdate="2003-01-01" firstname="Frank" gender="M" lastname="Kurmyshkin" nation="GER" license="300031" athleteid="6406">
              <ENTRIES>
                <ENTRY entrytime="00:09:07.65" entrycourse="LCM" eventid="2168" heatid="9616" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-01-19" name="Bayerische Meisterschaften lange Strecken" qualificationtime="00:09:19.65" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4441" nation="GER" region="02" clubid="6192" name="TSV Erding">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Sander" gender="M" lastname="Liebig" nation="GER" license="335431" athleteid="6193">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.35" entrycourse="SCM" eventid="1763" heatid="9380" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:10.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.47" entrycourse="SCM" eventid="1806" heatid="9419" lane="3">
                  <MEETINFO city="Erding" course="SCM" date="2019-10-05" name="4. Stadtwerke-Erding-Cup" qualificationtime="00:00:29.47" />
                </ENTRY>
                <ENTRY entrytime="00:02:22.87" entrycourse="SCM" eventid="1820" heatid="9430" lane="4">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:22.87" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.94" entrycourse="SCM" eventid="1834" heatid="9448" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:25.94" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.59" entrycourse="SCM" eventid="1985" heatid="9515" lane="6">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:31.59" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.53" entrycourse="SCM" eventid="2027" heatid="9543" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:04.53" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.32" entrycourse="SCM" eventid="2082" heatid="9570" lane="3">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-19" name="1. Internationaler Lechtal Cup" qualificationtime="00:02:36.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Andreas" gender="M" lastname="Rein" nation="GER" license="278278" athleteid="6201">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.00" entrycourse="SCM" eventid="1834" heatid="9451" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:23.05" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.98" entrycourse="SCM" eventid="1971" heatid="9495" lane="6">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:50.81" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.88" entrycourse="LCM" eventid="5307" heatid="9597" lane="6">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:25.88" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4452" nation="GER" region="02" clubid="6429" name="TSV Hohenbrunn-Riemerl.">
          <ATHLETES>
            <ATHLETE birthdate="2000-01-01" firstname="Adrien" gender="M" lastname="Cara" nation="GER" license="294598" athleteid="6430">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.72" entrycourse="LCM" eventid="1749" heatid="9363" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-03" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:01:51.72" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.29" entrycourse="SCM" eventid="1820" heatid="9433" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:05.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.00" entrycourse="SCM" eventid="1848" heatid="9469" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:02.00" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.29" entrycourse="SCM" eventid="1971" heatid="9495" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:52.29" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.39" entrycourse="SCM" eventid="2013" heatid="9537" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:57.86" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.44" entrycourse="LCM" eventid="2041" heatid="9559" lane="4">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:02:10.44" />
                </ENTRY>
                <ENTRY entrytime="00:04:04.73" entrycourse="LCM" eventid="2103" heatid="9613" lane="2">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:04:04.73" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Daniela" gender="F" lastname="Ernst" nation="GER" license="316890" athleteid="6438">
              <ENTRIES>
                <ENTRY entrytime="00:05:15.66" entrycourse="SCM" eventid="1771" heatid="9388" lane="1">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:05:15.66" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.32" entrycourse="SCM" eventid="1785" heatid="9401" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:04.32" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.60" entrycourse="SCM" eventid="1841" heatid="9460" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:00:31.15" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.48" entrycourse="SCM" eventid="2034" heatid="9553" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-06-01" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:30.69" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.85" entrycourse="SCM" eventid="2096" heatid="9606" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:19.85" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Alina" gender="F" lastname="Hermeking" nation="GER" license="290265" athleteid="6444">
              <ENTRIES>
                <ENTRY entrytime="00:02:34.15" entrycourse="SCM" eventid="2075" heatid="9564" lane="5">
                  <MEETINFO city="Bad Tölz" course="SCM" date="2019-02-24" name="DMS Bezirksdurchgang Oberbayern" qualificationtime="00:02:34.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:29.16" entrycourse="SCM" eventid="2096" heatid="9606" lane="1">
                  <MEETINFO city="Bad Tölz" course="SCM" date="2019-02-24" name="DMS Bezirksdurchgang Oberbayern" qualificationtime="00:02:29.16" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Sarah" gender="F" lastname="Hermeking" nation="GER" license="328767" athleteid="6447">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.38" entrycourse="SCM" eventid="1756" heatid="9372" lane="1">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:00:35.58" />
                </ENTRY>
                <ENTRY entrytime="00:02:48.59" entrycourse="SCM" eventid="1827" heatid="9438" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:51.10" />
                </ENTRY>
                <ENTRY entrytime="00:01:17.10" entrycourse="SCM" eventid="1992" heatid="9522" lane="5">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:18.65" />
                </ENTRY>
                <ENTRY entrytime="00:02:33.35" entrycourse="SCM" eventid="2075" heatid="9564" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:33.35" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Jette" gender="F" lastname="Lenz" nation="GER" license="348574" athleteid="6452">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.41" entrycourse="SCM" eventid="1059" heatid="9353" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-28" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:59.41" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.70" entrycourse="SCM" eventid="1799" heatid="9413" lane="1">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:09.70" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.64" entrycourse="SCM" eventid="1841" heatid="9460" lane="1">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:30.64" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.46" entrycourse="SCM" eventid="1978" heatid="9504" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:02:09.46" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.43" entrycourse="SCM" eventid="2034" heatid="9552" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:32.43" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.37" entrycourse="SCM" eventid="2089" heatid="9586" lane="5">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:27.37" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Carolin" gender="F" lastname="Seeger" nation="GER" license="311578" athleteid="6459">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.73" entrycourse="SCM" eventid="1059" heatid="9351" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:01.73" />
                </ENTRY>
                <ENTRY entrytime="00:04:40.00" entrycourse="SCM" eventid="5320" heatid="9474" lane="3">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-19" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:04:40.15" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.07" entrycourse="SCM" eventid="1978" heatid="9505" lane="4">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-21" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:02:11.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.33" entrycourse="SCM" eventid="2089" heatid="9580" lane="6">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:00:29.36" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Mara" gender="F" lastname="Sokac" nation="GER" license="360312" athleteid="6464">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.21" entrycourse="SCM" eventid="1059" heatid="9353" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:00:58.21" />
                </ENTRY>
                <ENTRY entrytime="00:01:09.50" entrycourse="SCM" eventid="1799" heatid="9413" lane="5">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:01:12.10" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.96" entrycourse="SCM" eventid="1841" heatid="9462" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-29" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:28.96" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.20" entrycourse="SCM" eventid="2006" heatid="9530" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:01:05.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.49" entrycourse="SCM" eventid="2089" heatid="9588" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-31" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:26.49" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2001-01-01" firstname="Sina" gender="F" lastname="Wappenschmidt" nation="GER" license="269801" athleteid="6470">
              <ENTRIES>
                <ENTRY entrytime="00:04:58.90" entrycourse="SCM" eventid="1771" heatid="9388" lane="3">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:05:09.84" />
                </ENTRY>
                <ENTRY entrytime="00:04:30.55" entrycourse="LCM" eventid="5320" heatid="9475" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-02" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:04:34.21" />
                </ENTRY>
                <ENTRY entrytime="00:17:33.54" entrycourse="SCM" eventid="5318" heatid="9479" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:18:16.81" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.16" entrycourse="SCM" eventid="1978" heatid="9505" lane="3">
                  <MEETINFO city="Berlin" course="LCM" date="2019-08-03" name="131. Deutsche Meisterschaften Schwimmen" qualificationtime="00:02:09.16" />
                </ENTRY>
                <ENTRY entrytime="00:02:24.20" entrycourse="SCM" eventid="2075" heatid="9567" lane="4">
                  <MEETINFO city="Ingolstadt" course="SCM" date="2019-02-03" name="DMS Bayernliga" qualificationtime="00:02:25.63" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.50" eventid="5314" heatid="9483" lane="4">
                  <MEETINFO city="München Obergiesing" date="2019-03-23" name="OMP Frühjahrsdurchgang - Jugend" qualificationtime="00:02:17.25" />
                </ENTRY>
                <ENTRY entrytime="00:01:48.50" eventid="2224" heatid="9618" lane="4" />
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4492" nation="GER" region="02" clubid="6346" name="TSV Vaterstetten">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Christian" gender="M" lastname="Arzberger" nation="GER" license="290446" athleteid="6347">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.61" entrycourse="LCM" eventid="1749" heatid="9362" lane="6">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-07" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:02:06.70" />
                </ENTRY>
                <ENTRY entrytime="00:01:07.79" entrycourse="SCM" eventid="1763" heatid="9383" lane="5">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:07.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.03" entrycourse="SCM" eventid="1820" heatid="9433" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:16.03" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.14" entrycourse="SCM" eventid="1848" heatid="9469" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:19.89" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.55" entrycourse="SCM" eventid="1971" heatid="9493" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:55.33" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.93" entrycourse="SCM" eventid="1985" heatid="9513" lane="4">
                  <MEETINFO city="Berlin" course="LCM" date="2019-05-30" name="Deutsche Jahrgangsmeisterschaften" qualificationtime="00:00:31.55" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.19" entrycourse="SCM" eventid="2027" heatid="9544" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:01:04.19" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.92" entrycourse="SCM" eventid="2082" heatid="9573" lane="1">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:32.28" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1988-01-01" firstname="Raul" gender="M" lastname="Garcia Alcaraz" nation="GER" license="399450" athleteid="6356">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.37" entrycourse="SCM" eventid="1971" heatid="9492" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:55.03" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.62" entrycourse="SCM" eventid="2027" heatid="9544" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:02.62" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.93" entrycourse="SCM" eventid="5307" heatid="9596" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:26.81" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Marlen Seraphine" gender="F" lastname="Görlach" nation="GER" license="306532" athleteid="6360">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.77" entrycourse="SCM" eventid="1059" heatid="9349" lane="2">
                  <MEETINFO city="Würzburg" course="LCM" date="2019-07-20" name="Bayerische Jahrgangsmeisterschaften" qualificationtime="00:01:02.77" />
                </ENTRY>
                <ENTRY entrytime="00:05:34.57" entrycourse="SCM" eventid="1771" heatid="9387" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:05:34.57" />
                </ENTRY>
                <ENTRY entrytime="00:01:12.97" entrycourse="SCM" eventid="1799" heatid="9410" lane="6">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:12.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:37.53" entrycourse="SCM" eventid="2075" heatid="9563" lane="5">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:37.53" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.32" entrycourse="SCM" eventid="2089" heatid="9580" lane="1">
                  <MEETINFO city="Kaufering" course="SCM" date="2019-01-20" name="1. Internationaler Lechtal Cup" qualificationtime="00:00:29.32" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Moritz" gender="M" lastname="Jung" nation="GER" license="295289" athleteid="6366">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.23" entrycourse="SCM" eventid="1749" heatid="9362" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:03.20" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.51" entrycourse="SCM" eventid="1778" heatid="9391" lane="6">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:01.51" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.01" entrycourse="SCM" eventid="1834" heatid="9447" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:26.01" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Johanna" gender="F" lastname="Latzel" nation="GER" license="375698" athleteid="6370">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.91" entrycourse="SCM" eventid="1785" heatid="9399" lane="5">
                  <MEETINFO city="München Obergiesing" course="SCM" date="2019-03-23" name="OMP Frühjahrsdurchgang - Offen/Minis" qualificationtime="00:01:11.91" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1996-01-01" firstname="Dominik" gender="M" lastname="Liguori" nation="GER" license="180738" athleteid="6372">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.04" entrycourse="SCM" eventid="1749" heatid="9364" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:59.65" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.24" entrycourse="SCM" eventid="1806" heatid="9421" lane="3">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:27.38" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.09" entrycourse="SCM" eventid="1834" heatid="9452" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:24.09" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.60" entrycourse="SCM" eventid="1971" heatid="9496" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:52.31" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.11" entrycourse="SCM" eventid="2013" heatid="9538" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:58.71" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.08" entrycourse="SCM" eventid="5307" heatid="9596" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:27.04" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Melissa" gender="F" lastname="Lux" nation="GER" license="287019" athleteid="6379">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.66" entrycourse="SCM" eventid="1785" heatid="9398" lane="3">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:01:12.66" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.18" entrycourse="SCM" eventid="2034" heatid="9551" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:33.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1999-01-01" firstname="Julius" gender="M" lastname="Schmid" nation="GER" license="223352" athleteid="6382">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.50" entrycourse="SCM" eventid="1749" heatid="9365" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:01:56.50" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.24" entrycourse="SCM" eventid="1778" heatid="9392" lane="2">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:58.83" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.63" entrycourse="SCM" eventid="1820" heatid="9431" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:02:14.07" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.51" entrycourse="LCM" eventid="1834" heatid="9449" lane="2">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:25.54" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.13" entrycourse="SCM" eventid="1971" heatid="9496" lane="5">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:53.13" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.10" entrycourse="LCM" eventid="5307" heatid="9595" lane="3">
                  <MEETINFO city="Karlsruhe" course="LCM" date="2019-05-31" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:00:27.10" />
                </ENTRY>
                <ENTRY entrytime="00:04:13.84" entrycourse="SCM" eventid="2103" heatid="9613" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:04:14.25" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Adrian" gender="M" lastname="Schoondermark" nation="GER" license="351659" athleteid="6390">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.91" entrycourse="SCM" eventid="1749" heatid="9361" lane="3">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-01-12" name="34. Augsburger Zirbelnuss-Schwimmen" qualificationtime="00:02:04.91" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.13" entrycourse="SCM" eventid="1834" heatid="9447" lane="5">
                  <MEETINFO city="Freising" course="LCM" date="2019-06-29" name="Kreisjahrgangsmeisterschaften Kreis6" qualificationtime="00:00:26.13" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.92" entrycourse="SCM" eventid="1848" heatid="9466" lane="4">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:02:21.92" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.39" entrycourse="SCM" eventid="1971" heatid="9491" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-02-09" name="Kreisjahrgangsmeisterschaften K6 Obb." qualificationtime="00:00:56.39" />
                </ENTRY>
                <ENTRY entrytime="00:04:33.45" entrycourse="SCM" eventid="2103" heatid="9609" lane="3">
                  <MEETINFO city="Bayreuth" course="LCM" date="2019-04-06" name="Bay. Meisterschaften mit SMK für 11 Jährige" qualificationtime="00:04:33.45" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="1997-01-01" firstname="Melina" gender="F" lastname="Uhl" nation="GER" license="245415" athleteid="6396">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.61" entrycourse="SCM" eventid="2089" heatid="9583" lane="2">
                  <MEETINFO city="Bayreuth" course="SCM" date="2019-02-02" name="DMS bay. Landesliga Durchgang Bayreuth" qualificationtime="00:00:28.61" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2003-01-01" firstname="Valerie" gender="F" lastname="Wende" nation="GER" license="325391" athleteid="6398">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.01" entrycourse="SCM" eventid="1059" heatid="9350" lane="4">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-13" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:02.92" />
                </ENTRY>
                <ENTRY entrytime="00:01:13.70" entrycourse="SCM" eventid="1799" heatid="9409" lane="5">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:01:13.25" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.28" entrycourse="SCM" eventid="2089" heatid="9584" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-10-12" name="Oberbayerische Kurzbahnmeisterschaft" qualificationtime="00:00:28.05" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.30" eventid="5316" heatid="9480" lane="3">
                  <MEETINFO city="Karlsruhe" date="2019-05-31" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:01:56.26" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.21" eventid="2232" heatid="9620" lane="5">
                  <MEETINFO city="Karlsruhe" date="2019-05-31" name="51. DM d. Masters Kurze Strecken" qualificationtime="00:01:42.21" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.33" eventid="5303" heatid="9614" lane="2">
                  <MEETINFO city="München Obergiesing" date="2019-03-23" name="OMP Frühjahrsdurchgang - Offen/Minis" qualificationtime="00:02:07.18" />
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4502" nation="GER" region="02" clubid="6426" name="TSV Zirndorf">
          <ATHLETES>
            <ATHLETE birthdate="1987-01-01" firstname="Thomas" gender="M" lastname="Almer" nation="GER" license="229594" athleteid="6427">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.45" eventid="1971" heatid="9491" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4529" nation="GER" region="02" clubid="5695" name="Turnverein Münchberg">
          <ATHLETES>
            <ATHLETE birthdate="2002-01-01" firstname="Valentin" gender="M" lastname="Schmiedel" nation="GER" license="289162" athleteid="5696">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.35" entrycourse="SCM" eventid="1763" heatid="9382" lane="1">
                  <MEETINFO city="Pegnitz" course="SCM" date="2019-10-05" name="2. CabrioSol Cup" qualificationtime="00:01:08.87" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5107" nation="GER" region="02" clubid="6636" name="TV 1860 Immenstadt">
          <ATHLETES>
            <ATHLETE birthdate="1999-01-01" firstname="Marcus" gender="M" lastname="Joas" nation="GER" license="161806" athleteid="6637">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.60" entrycourse="SCM" eventid="1971" heatid="9491" lane="1">
                  <MEETINFO city="Kaufbeuren" course="SCM" date="2019-03-24" name="18. Internationaler Buron Cup" qualificationtime="00:00:56.46" />
                </ENTRY>
                <ENTRY entrytime="00:04:18.07" entrycourse="SCM" eventid="2103" heatid="9612" lane="5">
                  <MEETINFO city="Kaufbeuren" course="SCM" date="2019-03-24" name="18. Internationaler Buron Cup" qualificationtime="00:04:17.51" />
                </ENTRY>
                <ENTRY entrytime="00:09:04.50" entrycourse="SCM" eventid="2168" heatid="9617" lane="1">
                  <MEETINFO city="Bad Saulgau" course="SCM" date="2019-10-06" name="3. Int. Bad Saulgauer Langstreckencup" qualificationtime="00:09:04.50" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2002-01-01" firstname="Simon" gender="M" lastname="Joas" nation="GER" license="282570" athleteid="6641">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.00" entrycourse="SCM" eventid="1749" heatid="9360" lane="4">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Augsburg" qualificationtime="00:02:03.05" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.26" entrycourse="SCM" eventid="1820" heatid="9431" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:20.26" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.50" entrycourse="SCM" eventid="1834" heatid="9445" lane="2">
                  <MEETINFO city="Obergünzburg" course="SCM" date="2019-05-04" name="28. Obergünzburger Schwimmfest" qualificationtime="00:00:25.84" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.35" entrycourse="SCM" eventid="1848" heatid="9469" lane="6">
                  <MEETINFO city="Kaufbeuren" course="SCM" date="2019-03-23" name="18. Internationaler Buron Cup" qualificationtime="00:02:19.35" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.20" entrycourse="SCM" eventid="1971" heatid="9490" lane="1">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Augsburg" qualificationtime="00:00:57.20" />
                </ENTRY>
                <ENTRY entrytime="00:05:02.25" entrycourse="SCM" eventid="1999" heatid="9527" lane="2">
                  <MEETINFO city="Immenstadt" course="SCM" date="2019-10-12" name="33. Internationales Immenstädter Schwimmfest" qualificationtime="00:05:02.25" />
                </ENTRY>
                <ENTRY entrytime="00:04:26.00" entrycourse="SCM" eventid="2103" heatid="9611" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-02-03" name="DMS bay. Landesliga Durchgang Augsburg" qualificationtime="00:04:23.14" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6812" nation="GER" region="02" clubid="6338" name="TV Kempten">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Thimo" gender="M" lastname="Thorandt" nation="GER" license="356235" athleteid="6339">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.97" entrycourse="SCM" eventid="1763" heatid="9381" lane="6">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:09.97" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.90" entrycourse="SCM" eventid="1820" heatid="9431" lane="6">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-19" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:20.90" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.54" entrycourse="SCM" eventid="1985" heatid="9511" lane="4">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-28" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:32.56" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.26" entrycourse="SCM" eventid="2027" heatid="9543" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:01:05.85" />
                </ENTRY>
                <ENTRY entrytime="00:02:31.84" entrycourse="SCM" eventid="2082" heatid="9571" lane="5">
                  <MEETINFO city="Augsburg" course="SCM" date="2019-05-18" name="Bezirks-Jahrgangsmeisterschaften und Masters" qualificationtime="00:02:31.84" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.43" entrycourse="SCM" eventid="5307" heatid="9593" lane="1">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:00:28.43" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4639" nation="GER" region="02" clubid="5820" name="WSV Bad Tölz">
          <ATHLETES>
            <ATHLETE birthdate="2004-01-01" firstname="Valentina" gender="F" lastname="Proverbio" nation="GER" license="346174" athleteid="5821">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.37" entrycourse="SCM" eventid="1059" heatid="9353" lane="1">
                  <MEETINFO city="Bad Reichenhall" course="SCM" date="2019-01-26" name="8. Rupertusthermen - Pokal-Schwimmen" qualificationtime="00:01:01.32" />
                </ENTRY>
                <ENTRY entrytime="00:01:10.23" entrycourse="SCM" eventid="1785" heatid="9400" lane="2">
                  <MEETINFO city="Riemerling" course="SCM" date="2019-09-29" name="Hohenbrunner Herbstschwimmfest" qualificationtime="00:01:11.01" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.70" entrycourse="SCM" eventid="1841" heatid="9457" lane="2">
                  <MEETINFO city="Regensburg" course="LCM" date="2019-05-11" name="Int. arena Swim Meeting" qualificationtime="00:00:31.43" />
                </ENTRY>
                <ENTRY entrytime="00:02:15.40" entrycourse="LCM" eventid="1978" heatid="9503" lane="3">
                  <MEETINFO city="Graz-Eggenberg" course="LCM" date="2019-04-26" name="Int. Ströck ATUS Graz Trophy" qualificationtime="00:02:16.79" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.81" entrycourse="SCM" eventid="2034" heatid="9553" lane="2">
                  <MEETINFO city="Bad Tölz" course="SCM" date="2019-06-29" name="Kreisjahrgangsmeisterschaften K3 Obb" qualificationtime="00:00:32.12" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.56" entrycourse="SCM" eventid="2089" heatid="9587" lane="1">
                  <MEETINFO city="Holzkirchen" course="SCM" date="2019-02-09" name="Kreiskurzbahnmeisterschaften K3 Obb." qualificationtime="00:00:27.56" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1062" code="BAY" course="SCM" gender="M" name="M 02" type="MAXIMUM">
      <AGEGROUP agemax="17" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:23.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:59.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:21.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:28.60">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:38.90">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:09.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:26.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:34.50">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.40">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:24.90">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.70">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:09.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.60">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.40">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="5333" code="BAY" course="SCM" gender="M" name="M bis 03" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:24.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:59.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:23.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.60">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:38.40">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:26.80">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:14.90">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:13.10">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.90">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:06.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="5339" code="BAY" course="SCM" gender="M" name="M offen" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="18" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:17.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:16.20">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:27.50">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:32.70">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:04.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:25.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:24.10">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.90">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:19.10">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:58.80">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.60">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:04.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1068" code="BAY" course="SCM" gender="F" name="W 03" type="MAXIMUM">
      <AGEGROUP agemax="16" agemin="16" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:35.90">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:35.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:31.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.20">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:19.60">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:54.40">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:12.90">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:38.20">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:33.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:21.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:34.90">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.40">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1080" code="BAY" course="SCM" gender="F" name="W bis 04" type="MAXIMUM">
      <AGEGROUP agemax="15" agemin="1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:37.20">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:57.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:21.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:57.30">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:13.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:39.20">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:34.20">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:22.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:38.90">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:14.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1072" code="BAY" course="SCM" gender="F" name="W offen" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="17" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:31.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.90">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:30.70">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.40">
          <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:16.50">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:29.10">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:48.90">
          <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.50">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:35.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:32.90">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:19.10">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:29.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.20">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:11.80">
          <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
