<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SG Fürth" version="11.61084">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Fürth" name="43. Fürther Kinderschwimmen" course="SCM" deadline="2018-11-04" hostclub="SG Fürth" hostclub.url="http://www.sgfuerth.de" organizer="SG Fürth" organizer.url="http://www.sgfuerth.de" reservecount="2" startmethod="1" timing="AUTOMATIC" state="BY" nation="GER">
      <AGEDATE value="2019-11-09" type="YEAR" />
      <POOL name="Hallebad am Scherbsgraben" lanemin="1" lanemax="6" />
      <FACILITY city="Fürth" name="Hallebad am Scherbsgraben" nation="GER" state="BY" street="Scherbsgraben 15" zip="90765" />
      <POINTTABLE pointtableid="3011" name="FINA Point Scoring" version="2018" />
      <CONTACT city="Fürth" email="meldungen@sgfuerth.de" name="Matthias Fuchs" phone="09118101172" street="Lavendelweg 47" zip="90768" />
      <SESSIONS>
        <SESSION date="2019-11-09" daytime="08:30" endtime="11:27" number="1" officialmeeting="08:15" teamleadermeeting="08:15" warmupfrom="08:00" warmupuntil="08:45">
          <EVENTS>
            <EVENT eventid="5668" daytime="08:40" gender="M" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="103" name="25m Rückenbeine ohne Brett" stroke="UNKNOWN" code="25 Rub" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7651" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7652" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7653" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7654" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25618" daytime="08:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25619" daytime="08:45" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7691" daytime="09:05" gender="M" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="501" name="25m Kraulbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7692" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7693" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7694" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7695" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25632" daytime="09:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25633" daytime="09:05" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25634" daytime="09:05" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5678" daytime="08:50" gender="M" number="5" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7659" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7660" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7661" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7662" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25622" daytime="08:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25623" daytime="08:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25624" daytime="08:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25625" daytime="08:55" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7696" daytime="09:05" gender="F" number="8" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="501" name="25m Kraulbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7697" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7698" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7699" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7700" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25635" daytime="09:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25636" daytime="09:10" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25637" daytime="09:10" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25638" daytime="09:10" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7706" daytime="09:55" gender="F" number="14" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="502" name="25m Delphinbeine o. Brett" stroke="UNKNOWN" code="25 Dob" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7707" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7708" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7709" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7710" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25658" daytime="09:55" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5674" daytime="08:45" gender="F" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="103" name="25m Rückenbeine ohne Brett" stroke="UNKNOWN" code="25 Rub" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7655" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7656" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7657" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7658" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25620" daytime="08:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25621" daytime="08:45" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5686" daytime="09:30" gender="M" number="9" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="101" name="25m Brustbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7667" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7668" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7669" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7670" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25639" daytime="09:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25640" daytime="09:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25641" daytime="09:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25642" daytime="09:35" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5664" daytime="08:35" gender="F" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7647" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7648" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7649" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7650" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25612" daytime="08:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25613" daytime="08:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25614" daytime="08:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25615" daytime="08:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25616" daytime="08:40" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25617" daytime="08:40" number="6" order="6" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5682" daytime="08:55" gender="F" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7663" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7664" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7665" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7666" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25626" daytime="08:55" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25627" daytime="08:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25628" daytime="09:00" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25629" daytime="09:00" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25630" daytime="09:00" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25631" daytime="09:00" number="6" order="6" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5694" daytime="09:40" gender="M" number="11" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7675" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7676" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7677" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7678" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25647" daytime="09:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25648" daytime="09:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25649" daytime="09:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25650" daytime="09:45" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5690" daytime="09:35" gender="F" number="10" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="101" name="25m Brustbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7671" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7672" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7673" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7674" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25643" daytime="09:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25644" daytime="09:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25645" daytime="09:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25646" daytime="09:40" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5698" daytime="09:45" gender="F" number="12" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7679" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7680" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7681" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7682" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25651" daytime="09:45" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25652" daytime="09:45" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25653" daytime="09:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25654" daytime="09:50" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25655" daytime="09:50" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25656" daytime="09:50" number="6" order="6" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1053" daytime="08:30" gender="M" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7646" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="1055" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="1054" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="2915" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25607" daytime="08:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25608" daytime="08:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25609" daytime="08:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25610" daytime="08:35" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25611" daytime="08:35" number="5" order="5" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7701" daytime="09:50" gender="M" number="13" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="502" name="25m Delphinbeine o. Brett" stroke="UNKNOWN" code="25 Dob" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7702" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7703" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7704" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7705" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25657" daytime="09:50" number="1" order="1" status="SEEDED" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2019-11-09" daytime="11:30" number="2" officialmeeting="11:00" teamleadermeeting="11:00" warmupfrom="10:30" warmupuntil="11:25">
          <EVENTS>
            <EVENT eventid="7773" daytime="15:15" gender="M" number="27" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7781" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7782" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7783" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7784" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7785" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7786" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7787" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25778" daytime="15:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25779" daytime="15:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25780" daytime="15:20" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25781" daytime="15:20" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25782" daytime="15:25" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25783" daytime="15:25" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25784" daytime="15:30" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5744" daytime="14:55" gender="F" number="26" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23817" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23818" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23819" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23820" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23821" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23822" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23823" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25761" daytime="14:55" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25762" daytime="15:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25763" daytime="15:00" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25764" daytime="15:00" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25765" daytime="15:00" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25766" daytime="15:05" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25767" daytime="15:05" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25768" daytime="15:05" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25769" daytime="15:05" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25770" daytime="15:05" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25771" daytime="15:10" number="11" order="11" status="SEEDED" />
                <HEAT heatid="25772" daytime="15:10" number="12" order="12" status="SEEDED" />
                <HEAT heatid="25773" daytime="15:10" number="13" order="13" status="SEEDED" />
                <HEAT heatid="25774" daytime="15:10" number="14" order="14" status="SEEDED" />
                <HEAT heatid="25775" daytime="15:10" number="15" order="15" status="SEEDED" />
                <HEAT heatid="25776" daytime="15:15" number="16" order="16" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7809" daytime="16:25" gender="F" number="30" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7818" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7819" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7820" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7821" agemax="11" agemin="11" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25798" daytime="16:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25799" daytime="16:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25800" daytime="16:25" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25801" daytime="16:25" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25802" daytime="16:25" number="5" order="5" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="13:00" gender="M" number="19" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7721" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1105" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1104" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1107" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1106" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1109" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25699" daytime="13:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25700" daytime="13:00" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7788" daytime="15:30" gender="F" number="28" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7789" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7790" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7791" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7792" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7793" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7794" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7795" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25785" daytime="15:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25786" daytime="15:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25787" daytime="15:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25788" daytime="15:35" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25789" daytime="15:40" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25790" daytime="15:40" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25791" daytime="15:45" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25792" daytime="15:45" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25793" daytime="15:45" number="9" order="9" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="16:50" gender="F" number="34" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7837" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7838" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7839" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7840" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7841" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7842" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7843" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25820" daytime="16:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25821" daytime="16:55" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25822" daytime="16:55" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25823" daytime="16:55" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25824" daytime="17:00" number="5" order="5" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5702" daytime="12:25" gender="M" number="17" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23782" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23783" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23784" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23785" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23786" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23787" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23788" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25673" daytime="12:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25674" daytime="12:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25675" daytime="12:30" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25676" daytime="12:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25677" daytime="12:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25678" daytime="12:30" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25679" daytime="12:35" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25680" daytime="12:35" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25681" daytime="12:35" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25682" daytime="12:35" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25683" daytime="12:40" number="11" order="11" status="SEEDED" />
                <HEAT heatid="25684" daytime="12:40" number="12" order="12" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5655" daytime="17:50" gender="M" number="37" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7870" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7871" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7872" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7873" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7874" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7875" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25848" daytime="17:50" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25849" daytime="17:50" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1177" daytime="11:30" gender="M" number="15" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7746" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7747" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7748" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7749" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7750" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7751" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25659" daytime="11:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25660" daytime="11:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25661" daytime="11:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25662" daytime="11:45" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25663" daytime="11:45" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25664" daytime="11:50" number="6" order="6" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5724" daytime="13:10" gender="M" number="21" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23796" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23797" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23798" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23799" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23800" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23801" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23802" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25704" daytime="13:10" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25705" daytime="13:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25706" daytime="13:15" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25707" daytime="13:15" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25708" daytime="13:15" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25709" daytime="13:20" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25710" daytime="13:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25711" daytime="13:20" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25712" daytime="13:20" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25713" daytime="13:25" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25714" daytime="13:25" number="11" order="11" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="17:25" gender="F" number="36" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7863" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7864" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7865" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7866" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7867" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7868" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7869" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25836" daytime="17:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25837" daytime="17:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25838" daytime="17:30" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25839" daytime="17:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25840" daytime="17:35" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25841" daytime="17:35" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25842" daytime="17:35" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25843" daytime="17:40" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25844" daytime="17:40" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25845" daytime="17:40" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25846" daytime="17:45" number="11" order="11" status="SEEDED" />
                <HEAT heatid="25847" daytime="17:45" number="12" order="12" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5740" daytime="14:40" gender="M" number="25" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23810" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23811" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23812" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23813" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23814" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23815" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23816" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25746" daytime="14:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25747" daytime="14:40" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25748" daytime="14:40" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25749" daytime="14:45" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25750" daytime="14:45" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25751" daytime="14:45" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25752" daytime="14:45" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25753" daytime="14:50" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25754" daytime="14:50" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25755" daytime="14:50" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25756" daytime="14:50" number="11" order="11" status="SEEDED" />
                <HEAT heatid="25757" daytime="14:50" number="12" order="12" status="SEEDED" />
                <HEAT heatid="25758" daytime="14:55" number="13" order="13" status="SEEDED" />
                <HEAT heatid="25759" daytime="14:55" number="14" order="14" status="SEEDED" />
                <HEAT heatid="25760" daytime="14:55" number="15" order="15" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5661" daytime="17:55" gender="F" number="38" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7876" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7877" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7878" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7879" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7880" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7881" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25850" daytime="17:55" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25851" daytime="18:00" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7804" daytime="16:20" gender="M" number="29" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7814" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7815" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7816" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7817" agemax="11" agemin="11" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25794" daytime="16:20" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25795" daytime="16:20" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25796" daytime="16:20" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25797" daytime="16:20" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5712" daytime="12:40" gender="F" number="18" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23789" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23790" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23791" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23792" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23793" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23794" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23795" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25685" daytime="12:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25686" daytime="12:45" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25687" daytime="12:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25688" daytime="12:45" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25689" daytime="12:45" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25690" daytime="12:50" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25691" daytime="12:50" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25692" daytime="12:50" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25693" daytime="12:55" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25694" daytime="12:55" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25695" daytime="12:55" number="11" order="11" status="SEEDED" />
                <HEAT heatid="25696" daytime="12:55" number="12" order="12" status="SEEDED" />
                <HEAT heatid="25697" daytime="12:55" number="13" order="13" status="SEEDED" />
                <HEAT heatid="25698" daytime="13:00" number="14" order="14" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" daytime="13:40" gender="M" number="23" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7759" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7760" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7761" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7762" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7763" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7764" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7765" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25729" daytime="13:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25730" daytime="14:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25731" daytime="14:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25732" daytime="14:05" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25733" daytime="14:10" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25734" daytime="14:10" number="6" order="6" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5728" daytime="13:25" gender="F" number="22" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23803" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23804" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23805" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23806" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23807" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23808" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23809" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25715" daytime="13:25" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25716" daytime="13:25" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25717" daytime="13:30" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25718" daytime="13:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25719" daytime="13:30" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25720" daytime="13:35" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25721" daytime="13:35" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25722" daytime="13:35" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25723" daytime="13:35" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25724" daytime="13:40" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25725" daytime="13:40" number="11" order="11" status="SEEDED" />
                <HEAT heatid="25726" daytime="13:40" number="12" order="12" status="SEEDED" />
                <HEAT heatid="25727" daytime="13:40" number="13" order="13" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="11:55" gender="F" number="16" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7753" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7754" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7755" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7756" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7757" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7758" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25665" daytime="11:55" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25666" daytime="12:00" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25667" daytime="12:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25668" daytime="12:05" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25669" daytime="12:10" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25670" daytime="12:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25671" daytime="12:20" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25672" daytime="12:20" number="8" order="8" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1189" daytime="17:00" gender="M" number="35" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7856" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7857" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7858" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7859" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7860" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7861" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7862" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25825" daytime="17:00" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25826" daytime="17:05" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25827" daytime="17:05" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25828" daytime="17:10" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25829" daytime="17:10" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25830" daytime="17:15" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25831" daytime="17:15" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25832" daytime="17:15" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25833" daytime="17:20" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25834" daytime="17:20" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25835" daytime="17:20" number="11" order="11" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="13:05" gender="F" number="20" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7722" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1112" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1113" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1114" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1115" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1116" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25701" daytime="13:05" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25702" daytime="13:05" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25703" daytime="13:10" number="3" order="3" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="14:15" gender="F" number="24" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7766" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7767" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7768" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7769" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7770" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7771" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7772" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25735" daytime="14:15" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25736" daytime="14:15" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25737" daytime="14:20" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25738" daytime="14:20" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25739" daytime="14:25" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25740" daytime="14:25" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25741" daytime="14:30" number="7" order="7" status="SEEDED" />
                <HEAT heatid="25742" daytime="14:30" number="8" order="8" status="SEEDED" />
                <HEAT heatid="25743" daytime="14:30" number="9" order="9" status="SEEDED" />
                <HEAT heatid="25744" daytime="14:35" number="10" order="10" status="SEEDED" />
                <HEAT heatid="25745" daytime="14:35" number="11" order="11" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="16:40" gender="M" number="33" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7830" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7831" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7832" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7833" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7834" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7835" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7836" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25816" daytime="16:40" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25817" daytime="16:45" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25818" daytime="16:45" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25819" daytime="16:50" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" daytime="16:30" gender="M" number="31" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23824" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23825" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23826" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23827" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23828" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23829" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23830" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25804" daytime="16:30" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25805" daytime="16:30" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25806" daytime="16:30" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25807" daytime="16:30" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25808" daytime="16:35" number="5" order="5" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1123" daytime="16:35" gender="F" number="32" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23831" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23832" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23833" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23834" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23835" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23836" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23837" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25809" daytime="16:35" number="1" order="1" status="SEEDED" />
                <HEAT heatid="25810" daytime="16:35" number="2" order="2" status="SEEDED" />
                <HEAT heatid="25811" daytime="16:35" number="3" order="3" status="SEEDED" />
                <HEAT heatid="25812" daytime="16:40" number="4" order="4" status="SEEDED" />
                <HEAT heatid="25813" daytime="16:40" number="5" order="5" status="SEEDED" />
                <HEAT heatid="25814" daytime="16:40" number="6" order="6" status="SEEDED" />
                <HEAT heatid="25815" daytime="16:40" number="7" order="7" status="SEEDED" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="4224" nation="GER" region="02" clubid="23845" name="Delphin 77 Herzogenaurach">
          <ATHLETES>
            <ATHLETE birthdate="2007-01-01" firstname="Fiona" gender="F" lastname="Baumann" nation="GER" license="403954" athleteid="23846">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.62" eventid="5712" heatid="25692" lane="5" />
                <ENTRY entrytime="00:00:49.42" eventid="5728" heatid="25723" lane="1" />
                <ENTRY entrytime="00:00:39.17" eventid="5744" heatid="25773" lane="2" />
                <ENTRY entrytime="00:01:44.65" eventid="7788" heatid="25790" lane="4" />
                <ENTRY entrytime="00:00:49.02" eventid="1123" heatid="25812" lane="2" />
                <ENTRY entrytime="00:01:27.66" eventid="1195" heatid="25845" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Amelie" gender="F" lastname="Bierlmeier" nation="GER" license="426838" athleteid="23853">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.13" eventid="5712" heatid="25691" lane="3" />
                <ENTRY entrytime="00:01:01.51" eventid="5728" heatid="25717" lane="3" />
                <ENTRY entrytime="00:00:55.21" eventid="5744" heatid="25764" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lena" gender="F" lastname="Bohrer" nation="GER" license="403950" athleteid="23857">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.35" eventid="5712" heatid="25695" lane="5" />
                <ENTRY entrytime="00:00:58.95" eventid="5728" heatid="25720" lane="5" />
                <ENTRY entrytime="00:01:58.13" eventid="1135" heatid="25739" lane="4" />
                <ENTRY entrytime="00:00:48.74" eventid="5744" heatid="25768" lane="1" />
                <ENTRY entrytime="00:00:58.76" eventid="1123" heatid="25809" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Theresa" gender="F" lastname="Dellermann" nation="GER" license="410601" athleteid="23863">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.06" eventid="5712" heatid="25697" lane="3" />
                <ENTRY entrytime="00:00:44.30" eventid="5728" heatid="25726" lane="4" />
                <ENTRY entrytime="00:01:43.26" eventid="1135" heatid="25744" lane="6" />
                <ENTRY entrytime="00:00:43.23" eventid="5744" heatid="25770" lane="4" />
                <ENTRY entrytime="00:01:45.00" eventid="7788" heatid="25790" lane="1" />
                <ENTRY entrytime="00:01:10.00" eventid="1123" heatid="25809" lane="1" />
                <ENTRY entrytime="00:01:28.36" eventid="1195" heatid="25844" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Andrea Jasmin" gender="F" lastname="Erm" nation="GER" license="999999" athleteid="23871">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5712" heatid="25688" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25719" lane="5" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="25765" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lene" gender="F" lastname="Friedrich" nation="GER" license="410600" athleteid="23875">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.51" eventid="5712" heatid="25698" lane="6" />
                <ENTRY entrytime="00:00:48.50" eventid="5728" heatid="25723" lane="4" />
                <ENTRY entrytime="00:00:37.49" eventid="5744" heatid="25775" lane="1" />
                <ENTRY entrytime="00:01:45.00" eventid="7788" heatid="25790" lane="5" />
                <ENTRY entrytime="00:01:28.40" eventid="1195" heatid="25844" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Thomas" gender="M" lastname="Hahn" nation="GER" license="999999" athleteid="23881">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5724" heatid="25704" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="25748" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Philipp" gender="M" lastname="Hardt" nation="GER" license="417042" athleteid="23884">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.19" eventid="5702" heatid="25683" lane="4" />
                <ENTRY entrytime="00:01:46.06" eventid="1141" heatid="25733" lane="6" />
                <ENTRY entrytime="00:00:37.04" eventid="5740" heatid="25758" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Simon" gender="M" lastname="Kamenik" nation="GER" license="410599" athleteid="23888">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.97" eventid="5702" heatid="25682" lane="3" />
                <ENTRY entrytime="00:00:46.40" eventid="5740" heatid="25752" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Mateo" gender="M" lastname="Kaufmair" nation="GER" license="382063" athleteid="23891">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.93" eventid="5702" heatid="25682" lane="6" />
                <ENTRY entrytime="00:00:49.19" eventid="5724" heatid="25711" lane="2" />
                <ENTRY entrytime="00:00:40.74" eventid="5740" heatid="25755" lane="3" />
                <ENTRY entrytime="00:01:44.28" eventid="7773" heatid="25781" lane="4" />
                <ENTRY entrytime="00:00:52.51" eventid="1117" heatid="25805" lane="3" />
                <ENTRY entrytime="00:01:27.37" eventid="1189" heatid="25832" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Luci" gender="F" lastname="Kitschke" nation="GER" license="417040" athleteid="23898">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.06" eventid="5712" heatid="25695" lane="2" />
                <ENTRY entrytime="00:00:50.72" eventid="5728" heatid="25722" lane="4" />
                <ENTRY entrytime="00:00:41.04" eventid="5744" heatid="25771" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Wilhelm" gender="M" lastname="Ruß" nation="GER" license="046841" athleteid="23902">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.81" eventid="5702" heatid="25680" lane="4" />
                <ENTRY entrytime="00:00:54.22" eventid="5724" heatid="25709" lane="5" />
                <ENTRY entrytime="00:01:57.00" eventid="1141" heatid="25731" lane="5" />
                <ENTRY entrytime="00:00:43.48" eventid="5740" heatid="25754" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="David" gender="M" lastname="Seefried" nation="GER" license="403947" athleteid="23907">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.67" eventid="5702" heatid="25680" lane="3" />
                <ENTRY entrytime="00:00:57.81" eventid="5724" heatid="25708" lane="1" />
                <ENTRY entrytime="00:00:45.34" eventid="5740" heatid="25753" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Jonathan" gender="M" lastname="Sopp" nation="GER" license="410602" athleteid="23911">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.51" eventid="5702" heatid="25679" lane="6" />
                <ENTRY entrytime="00:00:56.83" eventid="5724" heatid="25708" lane="4" />
                <ENTRY entrytime="00:01:57.00" eventid="1141" heatid="25731" lane="2" />
                <ENTRY entrytime="00:00:44.14" eventid="5740" heatid="25753" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emilja" gender="F" lastname="Stukelj" nation="GER" license="999999" athleteid="23916">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5712" heatid="25688" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25719" lane="2" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="25764" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Nilaksh Vikalp" gender="M" lastname="Yadav" nation="GER" license="046836" athleteid="23920">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="5702" heatid="25679" lane="4" />
                <ENTRY entrytime="00:00:54.85" eventid="5724" heatid="25709" lane="1" />
                <ENTRY entrytime="00:00:46.07" eventid="5740" heatid="25752" lane="4" />
                <ENTRY entrytime="00:01:37.00" eventid="1189" heatid="25829" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Paul" gender="M" lastname="Zitzmann" nation="GER" license="403945" athleteid="23925">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.86" eventid="5702" heatid="25680" lane="2" />
                <ENTRY entrytime="00:00:53.73" eventid="5724" heatid="25709" lane="3" />
                <ENTRY entrytime="00:00:41.66" eventid="5740" heatid="25755" lane="1" />
                <ENTRY entrytime="00:01:45.00" eventid="7773" heatid="25781" lane="5" />
                <ENTRY entrytime="00:01:35.24" eventid="1189" heatid="25830" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4271" nation="GER" region="02" clubid="24820" name="Post-SV Nürnberg">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Tobias" gender="M" lastname="Bonn" nation="GER" license="383469" athleteid="24821">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.40" eventid="5702" heatid="25684" lane="6" />
                <ENTRY entrytime="00:01:35.98" eventid="1141" heatid="25733" lane="2" />
                <ENTRY entrytime="00:00:35.00" eventid="5740" heatid="25759" lane="1" />
                <ENTRY entrytime="00:00:48.01" eventid="1117" heatid="25807" lane="6" />
                <ENTRY entrytime="00:01:18.56" eventid="1189" heatid="25833" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Hasset" gender="F" lastname="Efrem" nation="GER" license="392225" athleteid="24827">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.67" eventid="1111" heatid="25702" lane="5" />
                <ENTRY entrytime="00:01:48.00" eventid="1135" heatid="25743" lane="1" />
                <ENTRY entrytime="00:01:33.51" eventid="1171" heatid="25823" lane="3" />
                <ENTRY entrytime="00:01:14.86" eventid="1195" heatid="25847" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Daniel" gender="M" lastname="Hadersbrunner" nation="GER" license="392488" athleteid="24832">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.75" eventid="5702" heatid="25682" lane="5" />
                <ENTRY entrytime="00:00:49.90" eventid="5724" heatid="25711" lane="6" />
                <ENTRY entrytime="00:00:40.36" eventid="5740" heatid="25756" lane="5" />
                <ENTRY entrytime="00:01:29.63" eventid="1189" heatid="25831" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Marco" gender="M" lastname="Hadersbrunner" nation="GER" license="392487" athleteid="24837">
              <ENTRIES>
                <ENTRY entrytime="00:03:03.68" eventid="1177" heatid="25662" lane="2" />
                <ENTRY entrytime="00:01:47.98" eventid="1141" heatid="25732" lane="4" />
                <ENTRY entrytime="00:00:43.79" eventid="1117" heatid="25807" lane="3" />
                <ENTRY entrytime="00:01:27.75" eventid="1189" heatid="25832" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Simon" gender="M" lastname="Hadersbrunner" nation="GER" license="383461" athleteid="24842">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.13" eventid="5702" heatid="25684" lane="5" />
                <ENTRY entrytime="00:01:23.18" eventid="1103" heatid="25700" lane="4" />
                <ENTRY entrytime="00:00:31.89" eventid="5740" heatid="25760" lane="1" />
                <ENTRY entrytime="00:00:35.75" eventid="1117" heatid="25808" lane="3" />
                <ENTRY entrytime="00:01:12.86" eventid="1189" heatid="25834" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Leonora" gender="F" lastname="Hartmann" nation="GER" license="423845" athleteid="24848">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.51" eventid="5712" heatid="25688" lane="6" />
                <ENTRY entrytime="00:02:15.00" eventid="1135" heatid="25736" lane="5" />
                <ENTRY entrytime="00:00:35.00" eventid="7809" heatid="25799" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Timea Viola" gender="F" lastname="Heim" nation="GER" license="426097" athleteid="24852">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.00" eventid="1111" heatid="25702" lane="2" />
                <ENTRY entrytime="00:00:39.91" eventid="5744" heatid="25772" lane="3" />
                <ENTRY entrytime="00:00:47.68" eventid="1123" heatid="25813" lane="6" />
                <ENTRY entrytime="00:01:33.29" eventid="1195" heatid="25842" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Marie" gender="F" lastname="Hoppen" nation="GER" license="423843" athleteid="24862">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.39" eventid="5712" heatid="25691" lane="1" />
                <ENTRY entrytime="00:00:59.57" eventid="5728" heatid="25720" lane="6" />
                <ENTRY entrytime="00:00:50.22" eventid="5744" heatid="25766" lane="1" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25801" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="David" gender="M" lastname="Höhne" nation="GER" license="423839" athleteid="24857">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.00" eventid="5702" heatid="25678" lane="6" />
                <ENTRY entrytime="00:00:59.00" eventid="5724" heatid="25707" lane="5" />
                <ENTRY entrytime="00:00:58.00" eventid="5740" heatid="25749" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="7804" heatid="25794" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Elmercy" gender="F" lastname="Lulseged" nation="GER" license="426098" athleteid="24867">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.73" eventid="5712" heatid="25691" lane="2" />
                <ENTRY entrytime="00:00:52.35" eventid="5728" heatid="25722" lane="1" />
                <ENTRY entrytime="00:00:45.17" eventid="5744" heatid="25769" lane="4" />
                <ENTRY entrytime="00:00:26.50" eventid="7809" heatid="25800" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Johannes" gender="M" lastname="Lulseged" nation="GER" license="0" athleteid="24872">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.00" eventid="1053" heatid="25611" lane="6" />
                <ENTRY entrytime="00:00:25.00" eventid="5678" heatid="25625" lane="1" />
                <ENTRY entrytime="00:00:35.00" eventid="5686" heatid="25642" lane="1" />
                <ENTRY entrytime="00:00:29.00" eventid="5694" heatid="25650" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Rebekah" gender="F" lastname="Lulseged" nation="GER" license="383476" athleteid="24877">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.38" eventid="1135" heatid="25742" lane="5" />
                <ENTRY entrytime="00:00:37.88" eventid="5744" heatid="25775" lane="6" />
                <ENTRY entrytime="00:00:45.92" eventid="1123" heatid="25814" lane="6" />
                <ENTRY entrytime="00:01:52.63" eventid="1171" heatid="25821" lane="2" />
                <ENTRY entrytime="00:01:24.97" eventid="1195" heatid="25845" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Meggy" gender="F" lastname="Messel" nation="GER" license="423846" athleteid="24883">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.03" eventid="5712" heatid="25695" lane="1" />
                <ENTRY entrytime="00:00:49.40" eventid="5728" heatid="25723" lane="5" />
                <ENTRY entrytime="00:00:41.12" eventid="5744" heatid="25771" lane="5" />
                <ENTRY entrytime="00:00:19.94" eventid="7809" heatid="25802" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Samvel" gender="M" lastname="Mkrtchyan" nation="GER" license="426095" athleteid="24888">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.94" eventid="5702" heatid="25678" lane="1" />
                <ENTRY entrytime="00:00:54.11" eventid="5724" heatid="25709" lane="2" />
                <ENTRY entrytime="00:00:45.56" eventid="5740" heatid="25753" lane="6" />
                <ENTRY entrytime="00:00:23.00" eventid="7804" heatid="25797" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Michelle" gender="F" lastname="Möbus" nation="GER" license="423840" athleteid="24893">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.13" eventid="5712" heatid="25692" lane="6" />
                <ENTRY entrytime="00:00:50.25" eventid="5728" heatid="25722" lane="3" />
                <ENTRY entrytime="00:00:43.32" eventid="5744" heatid="25770" lane="5" />
                <ENTRY entrytime="00:00:23.60" eventid="7809" heatid="25802" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Sarah" gender="F" lastname="Olalowo" nation="GER" license="383462" athleteid="24898">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.00" eventid="1111" heatid="25702" lane="4" />
                <ENTRY entrytime="00:01:25.51" eventid="1135" heatid="25745" lane="3" />
                <ENTRY entrytime="00:01:30.36" eventid="1171" heatid="25824" lane="1" />
                <ENTRY entrytime="00:01:18.50" eventid="1195" heatid="25847" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Nick" gender="M" lastname="Rein" nation="GER" license="416115" athleteid="24903">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.10" eventid="5702" heatid="25681" lane="5" />
                <ENTRY entrytime="00:00:49.60" eventid="5724" heatid="25711" lane="5" />
                <ENTRY entrytime="00:00:41.81" eventid="5740" heatid="25755" lane="6" />
                <ENTRY entrytime="00:00:22.50" eventid="7804" heatid="25797" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Oskar" gender="M" lastname="Sonnenschein" nation="GER" license="423842" athleteid="24908">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.00" eventid="5702" heatid="25678" lane="4" />
                <ENTRY entrytime="00:00:47.93" eventid="5724" heatid="25712" lane="2" />
                <ENTRY entrytime="00:00:42.28" eventid="5740" heatid="25754" lane="3" />
                <ENTRY entrytime="00:00:25.47" eventid="7804" heatid="25796" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Maximilian" gender="M" lastname="Tatár" nation="GER" license="412059" athleteid="24913">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.06" eventid="5702" heatid="25681" lane="2" />
                <ENTRY entrytime="00:00:53.25" eventid="5724" heatid="25710" lane="1" />
                <ENTRY entrytime="00:00:45.37" eventid="5740" heatid="25753" lane="1" />
                <ENTRY entrytime="00:00:25.00" eventid="7804" heatid="25796" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Mikhael" gender="M" lastname="Varazhbitau" nation="GER" license="0" athleteid="24918">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.00" eventid="1053" heatid="25611" lane="5" />
                <ENTRY entrytime="00:00:38.00" eventid="5678" heatid="25623" lane="4" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="25641" lane="1" />
                <ENTRY entrytime="00:00:39.00" eventid="5694" heatid="25648" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lara" gender="F" lastname="Vogeler" nation="GER" license="0" athleteid="24923">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.00" eventid="5664" heatid="25616" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="5682" heatid="25630" lane="1" />
                <ENTRY entrytime="00:00:33.00" eventid="5698" heatid="25655" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="7706" heatid="25658" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2015-01-01" firstname="Roman" gender="M" lastname="Vogeler" nation="GER" license="0" athleteid="24928">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1053" heatid="25608" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25639" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lukas" gender="M" lastname="Westphal" nation="GER" license="412060" athleteid="24931">
              <ENTRIES>
                <ENTRY entrytime="00:03:09.85" eventid="1177" heatid="25662" lane="5" />
                <ENTRY entrytime="00:00:48.00" eventid="5724" heatid="25712" lane="5" />
                <ENTRY entrytime="00:00:40.18" eventid="5740" heatid="25756" lane="2" />
                <ENTRY entrytime="00:01:32.55" eventid="1189" heatid="25830" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lars" gender="M" lastname="Willums" nation="GER" license="423841" athleteid="24936">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.76" eventid="5702" heatid="25678" lane="5" />
                <ENTRY entrytime="00:00:57.99" eventid="5724" heatid="25708" lane="6" />
                <ENTRY entrytime="00:00:48.22" eventid="5740" heatid="25752" lane="5" />
                <ENTRY entrytime="00:00:30.00" eventid="7804" heatid="25795" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Leni" gender="F" lastname="Willums" nation="GER" license="0" athleteid="24941">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="5664" heatid="25616" lane="1" />
                <ENTRY entrytime="00:00:45.00" eventid="7696" heatid="25637" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="25652" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6524" nation="GER" region="02" clubid="25355" name="SC Regensburg">
          <ATHLETES>
            <ATHLETE birthdate="2012-01-01" firstname="Maxim" gender="M" lastname="Belyaev" nation="GER" license="000000" athleteid="25356">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.20" eventid="1053" heatid="25608" lane="4" />
                <ENTRY entrytime="NT" eventid="5668" heatid="25618" lane="5" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25632" lane="1" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25639" lane="2" />
                <ENTRY entrytime="00:00:33.08" eventid="5694" heatid="25649" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Luis" gender="M" lastname="Ewald" nation="GER" license="000000" athleteid="25362">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25607" lane="2" />
                <ENTRY entrytime="NT" eventid="5668" heatid="25618" lane="3" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25622" lane="5" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25632" lane="5" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25647" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Emilie" gender="F" lastname="Gierl" nation="GER" license="000000" athleteid="25368">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5674" heatid="25621" lane="6" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25635" lane="6" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25643" lane="1" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25652" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Alexander" gender="M" lastname="Hutchinson Riquelme" nation="GER" license="000000" athleteid="25373">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25618" lane="2" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25647" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Elias" gender="M" lastname="Jost" nation="GER" license="000000" athleteid="25376">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.11" eventid="1053" heatid="25609" lane="2" />
                <ENTRY entrytime="00:00:41.98" eventid="5668" heatid="25619" lane="1" />
                <ENTRY entrytime="00:00:42.10" eventid="7691" heatid="25633" lane="4" />
                <ENTRY entrytime="00:00:56.61" eventid="5686" heatid="25640" lane="4" />
                <ENTRY entrytime="00:00:34.02" eventid="5694" heatid="25649" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Sophia" gender="F" lastname="Löw" nation="GER" license="000000" athleteid="25382">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5674" heatid="25621" lane="1" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25643" lane="4" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25652" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Klara" gender="F" lastname="Nagler" nation="GER" license="000000" athleteid="25386">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25613" lane="1" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25620" lane="2" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25635" lane="2" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25643" lane="5" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25651" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Justus" gender="M" lastname="Rakow" nation="GER" license="000000" athleteid="25392">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25618" lane="1" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25647" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Emilian" gender="M" lastname="Rauch" nation="GER" license="000000" athleteid="25395">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25618" lane="4" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25647" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Leon" gender="M" lastname="Rauscher" nation="GER" license="000000" athleteid="25398">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.15" eventid="5668" heatid="25619" lane="2" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25622" lane="4" />
                <ENTRY entrytime="00:00:33.50" eventid="7691" heatid="25634" lane="3" />
                <ENTRY entrytime="00:00:34.60" eventid="5694" heatid="25649" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Frida" gender="F" lastname="Rosenbaum" nation="GER" license="000000" athleteid="25403">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25612" lane="4" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25620" lane="3" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25643" lane="2" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25651" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Johanna" gender="F" lastname="Spitzner" nation="GER" license="000000" athleteid="25408">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.29" eventid="5674" heatid="25621" lane="2" />
                <ENTRY entrytime="00:00:46.94" eventid="7696" heatid="25637" lane="2" />
                <ENTRY entrytime="00:00:31.93" eventid="5698" heatid="25656" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Antoni" gender="M" lastname="Swietlik" nation="GER" license="000000" athleteid="25412">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.27" eventid="5668" heatid="25619" lane="5" />
                <ENTRY entrytime="00:00:45.98" eventid="7691" heatid="25633" lane="5" />
                <ENTRY entrytime="00:00:30.22" eventid="5694" heatid="25650" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Oskar" gender="M" lastname="Swietlik" nation="GER" license="000000" athleteid="25416">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.84" eventid="5668" heatid="25619" lane="6" />
                <ENTRY entrytime="00:00:36.70" eventid="7691" heatid="25634" lane="5" />
                <ENTRY entrytime="00:00:33.12" eventid="5694" heatid="25649" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Caspar-Julius" gender="M" lastname="Wilke" nation="GER" license="368701" athleteid="25420">
              <ENTRIES>
                <ENTRY entrytime="00:02:32.68" eventid="1177" heatid="25664" lane="5" />
                <ENTRY entrytime="00:00:41.25" eventid="5702" heatid="25684" lane="2" />
                <ENTRY entrytime="00:01:28.08" eventid="1141" heatid="25734" lane="1" />
                <ENTRY entrytime="00:00:34.25" eventid="5740" heatid="25759" lane="2" />
                <ENTRY entrytime="00:01:20.36" eventid="1165" heatid="25819" lane="2" />
                <ENTRY entrytime="00:01:09.67" eventid="1189" heatid="25835" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Amilia" gender="F" lastname="Winkler" nation="GER" license="000000" athleteid="25427">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5674" heatid="25620" lane="1" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25635" lane="5" />
                <ENTRY entrytime="00:00:46.26" eventid="5698" heatid="25653" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4383" nation="GER" region="02" clubid="25435" name="SC Uttenreuth">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="David" gender="M" lastname="Felkel" nation="GER" license="0" athleteid="25436">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5702" heatid="25677" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="25748" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Yi Lin" gender="F" lastname="Gao" nation="GER" license="0" athleteid="25439">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.00" eventid="5712" heatid="25686" lane="4" />
                <ENTRY entrytime="00:01:15.00" eventid="5744" heatid="25761" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Paul" gender="M" lastname="Glanz" nation="GER" license="0" athleteid="25442">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.00" eventid="1053" heatid="25611" lane="2" />
                <ENTRY entrytime="00:00:25.00" eventid="5678" heatid="25625" lane="5" />
                <ENTRY entrytime="00:00:30.00" eventid="5694" heatid="25650" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lina" gender="F" lastname="Lederer" nation="GER" license="0" athleteid="25449">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.00" eventid="5664" heatid="25617" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" heatid="25637" lane="1" />
                <ENTRY entrytime="00:00:35.00" eventid="5698" heatid="25655" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Anna" gender="F" lastname="Schröter" nation="GER" license="0" athleteid="25453">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="5664" heatid="25615" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="5682" heatid="25630" lane="6" />
                <ENTRY entrytime="00:00:40.00" eventid="5690" heatid="25645" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Klara" gender="F" lastname="Schröter" nation="GER" license="0" athleteid="25457">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="5664" heatid="25616" lane="6" />
                <ENTRY entrytime="00:00:35.00" eventid="5682" heatid="25629" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="5690" heatid="25645" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6777" nation="GER" region="02" clubid="24066" name="Schwimmclub Schwandorf">
          <ATHLETES>
            <ATHLETE birthdate="2012-01-01" firstname="Luca" gender="M" lastname="Daucher" nation="GER" license="404783" athleteid="24067">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.02" eventid="1053" heatid="25610" lane="4" />
                <ENTRY entrytime="00:00:28.82" eventid="5678" heatid="25625" lane="6" />
                <ENTRY entrytime="00:00:36.77" eventid="7691" heatid="25634" lane="1" />
                <ENTRY entrytime="00:00:31.80" eventid="5694" heatid="25649" lane="4" />
                <ENTRY entrytime="NT" eventid="7701" heatid="25657" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Carlotta" gender="F" lastname="Fleischmann" nation="GER" license="374674" athleteid="24073">
              <ENTRIES>
                <ENTRY entrytime="00:03:30.08" eventid="1183" heatid="25668" lane="5" />
                <ENTRY entrytime="00:00:49.26" eventid="5728" heatid="25723" lane="2" />
                <ENTRY entrytime="00:01:56.51" eventid="1135" heatid="25739" lane="3" />
                <ENTRY entrytime="00:01:45.08" eventid="7788" heatid="25790" lane="6" />
                <ENTRY entrytime="00:00:50.51" eventid="1123" heatid="25811" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lucie" gender="F" lastname="Gebele" nation="GER" license="405006" athleteid="24085">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.57" eventid="5712" heatid="25687" lane="4" />
                <ENTRY entrytime="00:01:15.55" eventid="5728" heatid="25715" lane="5" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25735" lane="4" />
                <ENTRY entrytime="00:01:09.03" eventid="5744" heatid="25762" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Helena" gender="F" lastname="Gäntzle" nation="GER" license="405005" athleteid="24079">
              <ENTRIES>
                <ENTRY entrytime="00:03:18.57" eventid="1183" heatid="25670" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1111" heatid="25702" lane="6" />
                <ENTRY entrytime="00:00:40.34" eventid="5744" heatid="25772" lane="6" />
                <ENTRY entrytime="00:01:44.40" eventid="7788" heatid="25790" lane="3" />
                <ENTRY entrytime="00:00:46.94" eventid="1123" heatid="25813" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Andreas" gender="M" lastname="Hiltl" nation="GER" license="371456" athleteid="24090">
              <ENTRIES>
                <ENTRY entrytime="00:04:12.62" eventid="1177" heatid="25659" lane="3" />
                <ENTRY entrytime="00:01:05.54" eventid="5702" heatid="25675" lane="6" />
                <ENTRY entrytime="00:01:00.48" eventid="5724" heatid="25706" lane="4" />
                <ENTRY entrytime="00:00:45.60" eventid="5740" heatid="25752" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Knerer" nation="GER" license="404785" athleteid="24095">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5674" heatid="25620" lane="4" />
                <ENTRY entrytime="00:00:31.86" eventid="5682" heatid="25630" lane="4" />
                <ENTRY entrytime="00:00:44.97" eventid="7696" heatid="25637" lane="3" />
                <ENTRY entrytime="00:00:36.75" eventid="5698" heatid="25655" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emma" gender="F" lastname="Köhn" nation="GER" license="418818" athleteid="24100">
              <ENTRIES>
                <ENTRY entrytime="00:03:43.16" eventid="1183" heatid="25666" lane="3" />
                <ENTRY entrytime="00:00:56.40" eventid="5712" heatid="25693" lane="2" />
                <ENTRY entrytime="00:00:42.23" eventid="5744" heatid="25770" lane="3" />
                <ENTRY entrytime="00:01:55.44" eventid="7788" heatid="25788" lane="1" />
                <ENTRY entrytime="00:00:57.29" eventid="1123" heatid="25810" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Abby" gender="F" lastname="Lukas" nation="GER" license="374673" athleteid="24106">
              <ENTRIES>
                <ENTRY entrytime="00:03:27.71" eventid="1183" heatid="25668" lane="4" />
                <ENTRY entrytime="00:02:15.00" eventid="1111" heatid="25701" lane="4" />
                <ENTRY entrytime="00:00:45.59" eventid="5744" heatid="25769" lane="2" />
                <ENTRY entrytime="00:02:01.46" eventid="7788" heatid="25787" lane="6" />
                <ENTRY entrytime="00:00:57.34" eventid="1123" heatid="25810" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Aleksei" gender="M" lastname="Malikoski" nation="GER" license="390306" athleteid="24112">
              <ENTRIES>
                <ENTRY entrytime="00:03:16.36" eventid="1177" heatid="25661" lane="4" />
                <ENTRY entrytime="00:00:49.75" eventid="5724" heatid="25711" lane="1" />
                <ENTRY entrytime="00:00:38.19" eventid="5740" heatid="25757" lane="2" />
                <ENTRY entrytime="00:00:55.24" eventid="1117" heatid="25805" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Eva" gender="F" lastname="Matthes" nation="GER" license="000000" athleteid="24117">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.41" eventid="5664" heatid="25615" lane="1" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25620" lane="5" />
                <ENTRY entrytime="00:00:37.55" eventid="5682" heatid="25629" lane="2" />
                <ENTRY entrytime="00:00:34.37" eventid="5690" heatid="25646" lane="5" />
                <ENTRY entrytime="00:00:42.56" eventid="5698" heatid="25654" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Ida" gender="F" lastname="Matthes" nation="GER" license="416783" athleteid="24123">
              <ENTRIES>
                <ENTRY entrytime="00:05:46.11" eventid="1183" heatid="25665" lane="1" />
                <ENTRY entrytime="00:00:59.53" eventid="5712" heatid="25691" lane="6" />
                <ENTRY entrytime="00:02:16.28" eventid="1135" heatid="25736" lane="1" />
                <ENTRY entrytime="00:00:54.36" eventid="5744" heatid="25765" lane="2" />
                <ENTRY entrytime="00:02:17.73" eventid="7788" heatid="25785" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Paulina" gender="F" lastname="Plößl" nation="GER" license="374754" athleteid="24129">
              <ENTRIES>
                <ENTRY entrytime="00:04:10.70" eventid="1183" heatid="25665" lane="2" />
                <ENTRY entrytime="00:00:58.52" eventid="5712" heatid="25691" lane="4" />
                <ENTRY entrytime="00:02:06.48" eventid="1135" heatid="25737" lane="1" />
                <ENTRY entrytime="00:02:16.88" eventid="7788" heatid="25785" lane="5" />
                <ENTRY entrytime="00:00:59.17" eventid="1123" heatid="25809" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Hanna" gender="F" lastname="Rieder" nation="GER" license="390308" athleteid="24135">
              <ENTRIES>
                <ENTRY entrytime="00:03:39.57" eventid="1183" heatid="25667" lane="5" />
                <ENTRY entrytime="00:02:20.00" eventid="1111" heatid="25701" lane="2" />
                <ENTRY entrytime="00:00:46.31" eventid="5744" heatid="25769" lane="1" />
                <ENTRY entrytime="00:02:02.10" eventid="7788" heatid="25786" lane="3" />
                <ENTRY entrytime="00:00:56.68" eventid="1123" heatid="25810" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Victoria" gender="F" lastname="Schmid" nation="GER" license="421993" athleteid="24141">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.75" eventid="5728" heatid="25715" lane="1" />
                <ENTRY entrytime="00:01:10.29" eventid="5744" heatid="25761" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leonie" gender="F" lastname="Seger" nation="GER" license="390311" athleteid="24144">
              <ENTRIES>
                <ENTRY entrytime="00:03:18.65" eventid="1183" heatid="25670" lane="1" />
                <ENTRY entrytime="00:00:50.16" eventid="5728" heatid="25723" lane="6" />
                <ENTRY entrytime="00:00:40.11" eventid="5744" heatid="25772" lane="5" />
                <ENTRY entrytime="00:01:50.08" eventid="7788" heatid="25789" lane="6" />
                <ENTRY entrytime="00:00:50.68" eventid="1123" heatid="25811" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Zoe" gender="F" lastname="Seger" nation="GER" license="390312" athleteid="24150">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.30" eventid="5712" heatid="25696" lane="5" />
                <ENTRY entrytime="00:02:05.00" eventid="1135" heatid="25737" lane="4" />
                <ENTRY entrytime="00:00:43.25" eventid="5744" heatid="25770" lane="2" />
                <ENTRY entrytime="00:02:05.36" eventid="7788" heatid="25786" lane="5" />
                <ENTRY entrytime="00:00:48.60" eventid="1123" heatid="25812" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Anton" gender="M" lastname="Stiegler" nation="GER" license="421391" athleteid="24156">
              <ENTRIES>
                <ENTRY entrytime="00:01:22.69" eventid="5702" heatid="25673" lane="5" />
                <ENTRY entrytime="00:01:31.33" eventid="5724" heatid="25704" lane="5" />
                <ENTRY entrytime="00:01:38.51" eventid="5740" heatid="25746" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lara" gender="F" lastname="Wachtel" nation="GER" license="404786" athleteid="24160">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.50" eventid="5664" heatid="25617" lane="6" />
                <ENTRY entrytime="00:00:26.22" eventid="5682" heatid="25631" lane="1" />
                <ENTRY entrytime="00:00:47.95" eventid="5690" heatid="25645" lane="6" />
                <ENTRY entrytime="00:00:31.11" eventid="5698" heatid="25656" lane="1" />
                <ENTRY entrytime="NT" eventid="7706" heatid="25658" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Pauline" gender="F" lastname="Wiederer" nation="GER" license="390242" athleteid="24166">
              <ENTRIES>
                <ENTRY entrytime="00:03:53.12" eventid="1183" heatid="25666" lane="5" />
                <ENTRY entrytime="00:00:48.28" eventid="5728" heatid="25723" lane="3" />
                <ENTRY entrytime="00:02:05.54" eventid="1135" heatid="25737" lane="5" />
                <ENTRY entrytime="00:02:01.33" eventid="7788" heatid="25787" lane="1" />
                <ENTRY entrytime="00:00:54.49" eventid="1123" heatid="25811" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lina-Marie" gender="F" lastname="Zimmermann-Grünauer" nation="GER" license="420366" athleteid="24172">
              <ENTRIES>
                <ENTRY entrytime="00:04:11.21" eventid="1183" heatid="25665" lane="5" />
                <ENTRY entrytime="00:01:00.73" eventid="5712" heatid="25689" lane="3" />
                <ENTRY entrytime="00:02:10.32" eventid="1135" heatid="25736" lane="2" />
                <ENTRY entrytime="00:02:10.80" eventid="7788" heatid="25785" lane="4" />
                <ENTRY entrytime="00:01:03.81" eventid="1123" heatid="25809" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4302" nation="GER" region="02" clubid="24664" name="Schwimmfreunde Pegnitz">
          <ATHLETES>
            <ATHLETE birthdate="2008-01-01" firstname="Max" gender="M" lastname="Appelhans" nation="GER" license="382234" athleteid="24665">
              <ENTRIES>
                <ENTRY entrytime="00:03:16.75" eventid="1177" heatid="25661" lane="2" />
                <ENTRY entrytime="00:00:46.63" eventid="5724" heatid="25713" lane="5" />
                <ENTRY entrytime="00:00:38.77" eventid="5740" heatid="25756" lane="3" />
                <ENTRY entrytime="00:00:50.73" eventid="1117" heatid="25806" lane="1" />
                <ENTRY entrytime="00:01:29.14" eventid="1189" heatid="25831" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Hanna" gender="F" lastname="Büttner" nation="GER" license="419941" athleteid="24671">
              <ENTRIES>
                <ENTRY entrytime="00:03:30.45" eventid="1183" heatid="25668" lane="1" />
                <ENTRY entrytime="00:00:40.73" eventid="5728" heatid="25727" lane="5" />
                <ENTRY entrytime="00:01:31.23" eventid="1171" heatid="25824" lane="6" />
                <ENTRY entrytime="00:03:29.29" eventid="5661" heatid="25851" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jan" gender="M" lastname="Büttner" nation="GER" license="419943" athleteid="24676">
              <ENTRIES>
                <ENTRY entrytime="00:03:32.96" eventid="1177" heatid="25660" lane="4" />
                <ENTRY entrytime="00:00:46.80" eventid="5724" heatid="25713" lane="6" />
                <ENTRY entrytime="00:00:40.45" eventid="5740" heatid="25756" lane="1" />
                <ENTRY entrytime="00:01:48.00" eventid="7773" heatid="25781" lane="1" />
                <ENTRY entrytime="00:01:32.17" eventid="1189" heatid="25831" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Annika" gender="F" lastname="Reichel" nation="GER" license="419942" athleteid="24682">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.00" eventid="1183" heatid="25671" lane="2" />
                <ENTRY entrytime="00:00:46.65" eventid="5712" heatid="25698" lane="1" />
                <ENTRY entrytime="00:01:39.93" eventid="1135" heatid="25744" lane="4" />
                <ENTRY entrytime="00:03:29.82" eventid="5661" heatid="25851" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5147" nation="GER" region="02" clubid="23839" name="Schwimmgemeinschaft Fürth">
          <ATHLETES>
            <ATHLETE birthdate="2007-12-08" firstname="Philipp" gender="M" lastname="Adler" nation="GER" license="407267" athleteid="23977">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.87" entrycourse="SCM" eventid="5702" heatid="25676" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="7773" heatid="25778" lane="2" />
                <ENTRY entrytime="00:01:56.04" entrycourse="SCM" eventid="1189" heatid="25827" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Aidan" gender="M" lastname="Amelong" nation="GER" license="370804" athleteid="24492">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.74" eventid="5702" heatid="25682" lane="2" />
                <ENTRY entrytime="00:01:45.72" eventid="1141" heatid="25733" lane="1" />
                <ENTRY entrytime="00:01:18.54" eventid="1189" heatid="25833" lane="3" />
                <ENTRY entrytime="00:01:36.73" eventid="7773" heatid="25782" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Sina" gender="F" lastname="Amelong" nation="GER" license="378026" athleteid="24687">
              <ENTRIES>
                <ENTRY entrytime="00:03:23.58" eventid="1183" heatid="25669" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1111" heatid="25702" lane="1" />
                <ENTRY entrytime="00:01:05.80" eventid="7788" heatid="25793" lane="3" />
                <ENTRY entrytime="00:01:30.19" eventid="1195" heatid="25843" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sinan" gender="M" lastname="Arpert" nation="GER" license="297748" athleteid="24497">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.13" eventid="5702" heatid="25684" lane="4" />
                <ENTRY entrytime="00:01:27.19" eventid="1141" heatid="25734" lane="5" />
                <ENTRY entrytime="00:01:27.46" eventid="7773" heatid="25784" lane="6" />
                <ENTRY entrytime="00:03:02.69" eventid="5655" heatid="25849" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-03-07" firstname="Daniel" gender="M" lastname="Asev-Ajiyev" nation="GER" license="356304" athleteid="23981">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.81" entrycourse="SCM" eventid="5702" heatid="25680" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.35" entrycourse="SCM" eventid="5724" heatid="25708" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.82" entrycourse="SCM" eventid="5740" heatid="25753" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Marie" gender="F" lastname="Auerbach" nation="GER" license="391816" athleteid="24502">
              <ENTRIES>
                <ENTRY entrytime="00:01:47.35" eventid="1111" heatid="25703" lane="6" />
                <ENTRY entrytime="00:01:48.99" eventid="1135" heatid="25742" lane="3" />
                <ENTRY entrytime="00:01:39.94" eventid="7788" heatid="25791" lane="1" />
                <ENTRY entrytime="00:00:46.47" eventid="1123" heatid="25813" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Ida" gender="F" lastname="Baier" nation="GER" license="347848" athleteid="24945">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.96" eventid="5728" heatid="25725" lane="5" />
                <ENTRY entrytime="00:00:37.46" eventid="5744" heatid="25775" lane="5" />
                <ENTRY entrytime="00:00:39.92" eventid="1123" heatid="25815" lane="4" />
                <ENTRY entrytime="00:01:31.43" eventid="1195" heatid="25843" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lara" gender="F" lastname="Bamberger" nation="GER" license="362930" athleteid="24178">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.86" eventid="5712" heatid="25696" lane="4" />
                <ENTRY entrytime="00:00:47.65" eventid="5728" heatid="25724" lane="1" />
                <ENTRY entrytime="00:00:38.11" eventid="5744" heatid="25774" lane="5" />
                <ENTRY entrytime="00:00:50.74" eventid="1123" heatid="25811" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-23" firstname="Rebekka" gender="F" lastname="Behring" nation="GER" license="407272" athleteid="24482">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.00" eventid="5728" heatid="25717" lane="2" />
                <ENTRY entrytime="00:01:04.00" eventid="5744" heatid="25762" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Max Eric" gender="M" lastname="Besecke" nation="GER" license="406834" athleteid="24692">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1141" heatid="25730" lane="1" />
                <ENTRY entrytime="00:01:02.37" eventid="5740" heatid="25748" lane="6" />
                <ENTRY entrytime="00:02:05.00" eventid="1189" heatid="25826" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Alarice" gender="F" lastname="Bitz" nation="GER" athleteid="24696">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25612" lane="2" />
                <ENTRY entrytime="NT" eventid="5682" heatid="25626" lane="4" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25643" lane="6" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25652" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Benedek" gender="M" lastname="Boha" nation="GER" license="666666" athleteid="24701">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1177" heatid="25659" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="1141" heatid="25732" lane="6" />
                <ENTRY entrytime="NT" eventid="7773" heatid="25778" lane="4" />
                <ENTRY entrytime="00:01:40.00" eventid="1189" heatid="25829" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Dina" gender="F" lastname="Boha" nation="GER" license="391813" athleteid="24507">
              <ENTRIES>
                <ENTRY entrytime="00:02:47.51" eventid="1183" heatid="25672" lane="3" />
                <ENTRY entrytime="00:01:38.74" eventid="1135" heatid="25745" lane="6" />
                <ENTRY entrytime="00:01:30.09" eventid="7788" heatid="25793" lane="5" />
                <ENTRY entrytime="00:01:13.15" eventid="1195" heatid="25847" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-04-17" firstname="Daniel" gender="M" lastname="Bramigk" nation="GER" license="420770" athleteid="23990">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.48" entrycourse="SCM" eventid="5724" heatid="25707" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:48.64" entrycourse="SCM" eventid="5740" heatid="25752" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:44.78" entrycourse="LCM" eventid="1189" heatid="25829" lane="6">
                  <MEETINFO course="LCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Anastasia" gender="F" lastname="Chochlow" nation="GER" license="392745" athleteid="24706">
              <ENTRIES>
                <ENTRY entrytime="00:03:29.58" eventid="1183" heatid="25668" lane="2" />
                <ENTRY entrytime="00:00:02.00" eventid="1111" heatid="25703" lane="3" />
                <ENTRY entrytime="00:01:53.07" eventid="7788" heatid="25788" lane="2" />
                <ENTRY entrytime="00:01:35.19" eventid="1195" heatid="25841" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lena" gender="F" lastname="Clausen" nation="GER" license="420945" athleteid="24512">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.53" eventid="5712" heatid="25689" lane="6" />
                <ENTRY entrytime="00:01:04.27" eventid="5728" heatid="25717" lane="6" />
                <ENTRY entrytime="00:01:01.92" eventid="5744" heatid="25762" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="7809" heatid="25798" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Simon" gender="M" lastname="Clausen" nation="GER" athleteid="24517">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.38" eventid="1053" heatid="25609" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="7691" heatid="25633" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="5686" heatid="25640" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Helena" gender="F" lastname="Dautermann" nation="GER" license="393633" athleteid="24950">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.47" eventid="5712" heatid="25698" lane="2" />
                <ENTRY entrytime="00:00:46.68" eventid="5728" heatid="25724" lane="2" />
                <ENTRY entrytime="00:01:42.99" eventid="1135" heatid="25744" lane="1" />
                <ENTRY entrytime="00:00:38.99" eventid="5744" heatid="25774" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Simon" gender="M" lastname="Dieret" nation="GER" license="331161" athleteid="23840">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.62" eventid="5724" heatid="25714" lane="1" />
                <ENTRY entrytime="00:00:35.24" eventid="5740" heatid="25759" lane="6" />
                <ENTRY entrytime="00:01:33.75" eventid="7773" heatid="25783" lane="1" />
                <ENTRY entrytime="00:00:41.54" eventid="1117" heatid="25808" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Daniel" gender="M" lastname="Ehnis" nation="GER" license="378024" athleteid="24711">
              <ENTRIES>
                <ENTRY entrytime="00:03:57.93" eventid="1177" heatid="25660" lane="1" />
                <ENTRY entrytime="00:02:03.30" eventid="1141" heatid="25730" lane="2" />
                <ENTRY entrytime="00:02:06.48" eventid="7773" heatid="25779" lane="5" />
                <ENTRY entrytime="00:01:45.32" eventid="1189" heatid="25828" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Julia" gender="F" lastname="Ehnis" nation="GER" athleteid="24716">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.36" eventid="5664" heatid="25615" lane="4" />
                <ENTRY entrytime="00:00:48.60" eventid="5682" heatid="25628" lane="5" />
                <ENTRY entrytime="00:00:48.00" eventid="7696" heatid="25637" lane="5" />
                <ENTRY entrytime="00:00:45.51" eventid="5698" heatid="25654" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-02-15" firstname="Jakob" gender="M" lastname="Freund" nation="GER" license="331165" athleteid="23994">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.37" entrycourse="SCM" eventid="5702" heatid="25679" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.97" entrycourse="SCM" eventid="5724" heatid="25706" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.92" entrycourse="SCM" eventid="5740" heatid="25750" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:03.23" entrycourse="SCM" eventid="1117" heatid="25804" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Anna" gender="F" lastname="Fuchs" nation="GER" license="346281" athleteid="24955">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.85" eventid="5712" heatid="25697" lane="2" />
                <ENTRY entrytime="00:01:51.10" eventid="1135" heatid="25741" lane="4" />
                <ENTRY entrytime="00:00:39.66" eventid="5744" heatid="25773" lane="6" />
                <ENTRY entrytime="00:00:20.00" eventid="7809" heatid="25802" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lia Sophie" gender="F" lastname="Fuchs" nation="GER" license="420938" athleteid="24721">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.38" eventid="5664" heatid="25615" lane="5" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25621" lane="5" />
                <ENTRY entrytime="00:00:31.58" eventid="5682" heatid="25630" lane="3" />
                <ENTRY entrytime="00:00:33.75" eventid="5698" heatid="25655" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Maximilian" gender="M" lastname="Fuchs" nation="GER" license="342442" athleteid="24960">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.36" eventid="5702" heatid="25683" lane="3" />
                <ENTRY entrytime="00:01:35.51" eventid="1141" heatid="25733" lane="4" />
                <ENTRY entrytime="00:01:25.77" eventid="1189" heatid="25832" lane="3" />
                <ENTRY entrytime="00:00:37.07" eventid="5740" heatid="25758" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Linnea Emilia" gender="F" lastname="Glößinger" nation="GER" license="389377" athleteid="24726">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.84" eventid="5664" heatid="25616" lane="2" />
                <ENTRY entrytime="00:00:36.63" eventid="5682" heatid="25629" lane="4" />
                <ENTRY entrytime="00:00:00.50" eventid="5690" heatid="25646" lane="3" />
                <ENTRY entrytime="00:00:36.14" eventid="5698" heatid="25655" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Anton" gender="M" lastname="Grießinger" nation="GER" license="362946" athleteid="24521">
              <ENTRIES>
                <ENTRY entrytime="00:01:26.58" eventid="1103" heatid="25700" lane="2" />
                <ENTRY entrytime="00:01:40.44" eventid="1141" heatid="25733" lane="5" />
                <ENTRY entrytime="00:01:27.92" eventid="7773" heatid="25783" lane="4" />
                <ENTRY entrytime="00:01:12.39" eventid="1189" heatid="25835" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Leyan Su" gender="F" lastname="Gülec" nation="GER" license="377883" athleteid="24965">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.50" eventid="5728" heatid="25727" lane="2" />
                <ENTRY entrytime="00:00:34.78" eventid="5744" heatid="25776" lane="4" />
                <ENTRY entrytime="00:00:41.75" eventid="1123" heatid="25815" lane="5" />
                <ENTRY entrytime="00:01:20.17" eventid="1195" heatid="25846" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Annika" gender="F" lastname="Haas" nation="GER" license="555555" athleteid="24183">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25718" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Maria Magdalena" gender="F" lastname="Haußwald" nation="GER" athleteid="24970">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.14" eventid="5712" heatid="25693" lane="6" />
                <ENTRY entrytime="00:00:52.18" eventid="5728" heatid="25722" lane="5" />
                <ENTRY entrytime="00:00:44.39" eventid="5744" heatid="25770" lane="6" />
                <ENTRY entrytime="00:01:43.59" eventid="1195" heatid="25840" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lilith" gender="F" lastname="Heidenreich" nation="GER" license="420940" athleteid="24526">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.43" eventid="5712" heatid="25687" lane="1" />
                <ENTRY entrytime="00:01:05.81" eventid="5744" heatid="25762" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Louisa" gender="F" lastname="Heidenreich" nation="GER" license="420942" athleteid="24529">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.76" eventid="5664" heatid="25614" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="25653" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Lorena" gender="F" lastname="Heinl" nation="GER" license="407278" athleteid="24975">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.28" eventid="5712" heatid="25696" lane="2" />
                <ENTRY entrytime="00:01:48.00" eventid="1135" heatid="25743" lane="5" />
                <ENTRY entrytime="00:00:49.00" eventid="5744" heatid="25767" lane="2" />
                <ENTRY entrytime="00:00:58.00" eventid="5728" heatid="25720" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Luisa" gender="F" lastname="Heyert" nation="GER" license="347335" athleteid="24532">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.65" eventid="5712" heatid="25696" lane="3" />
                <ENTRY entrytime="00:00:42.56" eventid="5728" heatid="25727" lane="6" />
                <ENTRY entrytime="00:01:30.77" eventid="7788" heatid="25793" lane="6" />
                <ENTRY entrytime="00:01:20.37" eventid="1195" heatid="25846" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Tobias" gender="M" lastname="Heyert" nation="GER" license="306630" athleteid="24537">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.65" eventid="5724" heatid="25714" lane="3" />
                <ENTRY entrytime="00:00:29.85" eventid="5740" heatid="25760" lane="2" />
                <ENTRY entrytime="00:01:16.78" eventid="1165" heatid="25819" lane="4" />
                <ENTRY entrytime="00:02:49.82" eventid="5655" heatid="25849" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Alissa" gender="F" lastname="Hilz" nation="GER" athleteid="24731">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25685" lane="4" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25735" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Julianna" gender="F" lastname="Jahn" nation="GER" athleteid="24542">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5728" heatid="25716" lane="6" />
                <ENTRY entrytime="00:01:10.00" eventid="5744" heatid="25761" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Emil" gender="M" lastname="Jeske" nation="GER" license="378027" athleteid="24734">
              <ENTRIES>
                <ENTRY entrytime="00:03:02.16" eventid="1177" heatid="25662" lane="4" />
                <ENTRY entrytime="00:01:50.00" eventid="1103" heatid="25699" lane="1" />
                <ENTRY entrytime="00:01:33.44" eventid="1165" heatid="25818" lane="3" />
                <ENTRY entrytime="00:03:00.00" eventid="5655" heatid="25849" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Vanessa" gender="F" lastname="Kenner" nation="GER" license="362937" athleteid="24185">
              <ENTRIES>
                <ENTRY entrytime="00:03:50.34" eventid="1183" heatid="25666" lane="2" />
                <ENTRY entrytime="00:02:00.99" eventid="1171" heatid="25821" lane="6" />
                <ENTRY entrytime="00:04:45.00" eventid="5661" heatid="25850" lane="2" />
                <ENTRY entrytime="00:02:10.00" eventid="1111" heatid="25701" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Max" gender="M" lastname="Keyser" nation="GER" license="420769" athleteid="24190">
              <ENTRIES>
                <ENTRY entrytime="00:02:59.12" eventid="1177" heatid="25663" lane="5" />
                <ENTRY entrytime="00:01:40.00" eventid="1103" heatid="25700" lane="6" />
                <ENTRY entrytime="00:03:40.00" eventid="5655" heatid="25848" lane="2" />
                <ENTRY entrytime="00:00:33.21" eventid="5740" heatid="25759" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Timm" gender="M" lastname="Laus" nation="GER" license="362943" athleteid="24195">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.69" eventid="5702" heatid="25679" lane="1" />
                <ENTRY entrytime="00:00:55.63" eventid="5724" heatid="25708" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="7773" heatid="25779" lane="4" />
                <ENTRY entrytime="00:01:55.00" eventid="1165" heatid="25816" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Luca" gender="M" lastname="Lautenschlager" nation="GER" license="404302" athleteid="23931">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.06" eventid="1053" heatid="25610" lane="3" />
                <ENTRY entrytime="00:00:35.41" eventid="5678" heatid="25624" lane="6" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="25641" lane="4" />
                <ENTRY entrytime="00:00:39.64" eventid="5694" heatid="25648" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Nils" gender="M" lastname="Lautenschlager" nation="GER" license="372637" athleteid="23936">
              <ENTRIES>
                <ENTRY entrytime="00:02:15.00" eventid="1141" heatid="25729" lane="2" />
                <ENTRY entrytime="00:00:55.19" eventid="5724" heatid="25709" lane="6" />
                <ENTRY entrytime="00:00:27.00" eventid="7804" heatid="25796" lane="5" />
                <ENTRY entrytime="00:02:15.00" eventid="1189" heatid="25825" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Edwin" gender="M" lastname="Lichtenwald" nation="GER" athleteid="24739">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.31" eventid="1053" heatid="25609" lane="4" />
                <ENTRY entrytime="00:00:33.54" eventid="5678" heatid="25624" lane="2" />
                <ENTRY entrytime="00:00:00.50" eventid="5686" heatid="25642" lane="2" />
                <ENTRY entrytime="00:00:37.22" eventid="5694" heatid="25648" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Livia" gender="F" lastname="Lichtenwald" nation="GER" license="393386" athleteid="24744">
              <ENTRIES>
                <ENTRY entrytime="00:03:22.51" eventid="1183" heatid="25669" lane="2" />
                <ENTRY entrytime="00:01:48.78" eventid="1111" heatid="25702" lane="3" />
                <ENTRY entrytime="00:01:46.72" eventid="1135" heatid="25743" lane="2" />
                <ENTRY entrytime="00:01:31.33" eventid="1195" heatid="25843" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Finn" gender="M" lastname="Martin" nation="GER" license="355301" athleteid="24200">
              <ENTRIES>
                <ENTRY entrytime="00:03:01.34" eventid="1177" heatid="25663" lane="6" />
                <ENTRY entrytime="00:01:40.91" eventid="1103" heatid="25699" lane="3" />
                <ENTRY entrytime="00:00:33.03" eventid="5740" heatid="25760" lane="6" />
                <ENTRY entrytime="00:03:45.00" eventid="5655" heatid="25848" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ida" gender="F" lastname="Martin" nation="GER" license="362939" athleteid="24205">
              <ENTRIES>
                <ENTRY entrytime="00:03:36.02" eventid="1183" heatid="25667" lane="2" />
                <ENTRY entrytime="00:02:17.91" eventid="1135" heatid="25736" lane="6" />
                <ENTRY entrytime="00:00:55.59" eventid="1123" heatid="25810" lane="2" />
                <ENTRY entrytime="00:01:42.54" eventid="1195" heatid="25840" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lasse" gender="M" lastname="Martin" nation="GER" license="000000" athleteid="25466">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25607" lane="3" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25632" lane="2" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25647" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Cosima" gender="F" lastname="Nahr" nation="GER" license="376904" athleteid="23941">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.56" eventid="5728" heatid="25721" lane="3" />
                <ENTRY entrytime="00:01:58.57" eventid="1135" heatid="25739" lane="5" />
                <ENTRY entrytime="00:00:26.00" eventid="7809" heatid="25801" lane="6" />
                <ENTRY entrytime="00:02:10.00" eventid="1195" heatid="25836" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Julius" gender="M" lastname="Nahr" nation="GER" license="416999" athleteid="23946">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.06" eventid="1053" heatid="25608" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="7691" heatid="25633" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="25641" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Julia" gender="F" lastname="Okner" nation="GER" athleteid="23950">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.38" eventid="5712" heatid="25685" lane="3" />
                <ENTRY entrytime="00:01:30.12" eventid="5744" heatid="25761" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jonas" gender="M" lastname="Penz" nation="GER" license="392570" athleteid="24210">
              <ENTRIES>
                <ENTRY entrytime="00:04:00.43" eventid="1177" heatid="25660" lane="6" />
                <ENTRY entrytime="00:00:53.53" eventid="5724" heatid="25710" lane="6" />
                <ENTRY entrytime="00:00:41.53" eventid="5740" heatid="25755" lane="2" />
                <ENTRY entrytime="00:01:42.69" eventid="1189" heatid="25829" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lara" gender="F" lastname="Penz" nation="GER" license="362938" athleteid="24215">
              <ENTRIES>
                <ENTRY entrytime="00:03:26.58" eventid="1183" heatid="25668" lane="3" />
                <ENTRY entrytime="00:00:36.68" eventid="5744" heatid="25775" lane="3" />
                <ENTRY entrytime="00:00:44.22" eventid="1123" heatid="25814" lane="2" />
                <ENTRY entrytime="00:03:37.69" eventid="5661" heatid="25851" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-13" firstname="Laurenz" gender="M" lastname="Raum" nation="GER" license="392567" athleteid="24489">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.00" eventid="5702" heatid="25676" lane="1" />
                <ENTRY entrytime="00:00:59.00" eventid="5740" heatid="25749" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lian" gender="M" lastname="Richter" nation="GER" license="406841" athleteid="24749">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1141" heatid="25730" lane="5" />
                <ENTRY entrytime="00:00:29.15" eventid="7804" heatid="25796" lane="1" />
                <ENTRY entrytime="NT" eventid="1165" heatid="25816" lane="5" />
                <ENTRY entrytime="00:02:25.28" eventid="1189" heatid="25825" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lisa" gender="F" lastname="Rischbeck" nation="GER" license="666666" athleteid="24754">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1135" heatid="25737" lane="2" />
                <ENTRY entrytime="NT" eventid="7788" heatid="25785" lane="6" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25798" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1195" heatid="25837" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Theo" gender="M" lastname="Rischbeck" nation="GER" license="666666" athleteid="24759">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.19" eventid="1053" heatid="25610" lane="5" />
                <ENTRY entrytime="00:00:33.82" eventid="5678" heatid="25624" lane="5" />
                <ENTRY entrytime="00:00:00.45" eventid="5686" heatid="25642" lane="4" />
                <ENTRY entrytime="00:00:36.23" eventid="5694" heatid="25648" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ronja" gender="F" lastname="Rosenthal" nation="GER" license="389376" athleteid="24764">
              <ENTRIES>
                <ENTRY entrytime="00:03:57.10" eventid="1183" heatid="25666" lane="6" />
                <ENTRY entrytime="00:01:49.69" eventid="1135" heatid="25742" lane="1" />
                <ENTRY entrytime="00:01:39.75" eventid="1171" heatid="25823" lane="5" />
                <ENTRY entrytime="00:01:32.28" eventid="1195" heatid="25842" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Leana Isabel" gender="F" lastname="Rother" nation="GER" license="379366" athleteid="23953">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.56" eventid="5728" heatid="25721" lane="4" />
                <ENTRY entrytime="00:01:58.44" eventid="1135" heatid="25739" lane="2" />
                <ENTRY entrytime="00:00:26.00" eventid="7809" heatid="25801" lane="1" />
                <ENTRY entrytime="00:01:53.91" eventid="1195" heatid="25839" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Theo" gender="M" lastname="Rother" nation="GER" athleteid="24769">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.25" eventid="1053" heatid="25610" lane="2" />
                <ENTRY entrytime="00:00:29.52" eventid="5678" heatid="25624" lane="3" />
                <ENTRY entrytime="00:00:00.45" eventid="5686" heatid="25642" lane="3" />
                <ENTRY entrytime="00:00:31.79" eventid="5694" heatid="25649" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Timon Sebastian" gender="M" lastname="Rother" nation="GER" license="406840" athleteid="23958">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.19" eventid="1053" heatid="25610" lane="1" />
                <ENTRY entrytime="00:00:35.43" eventid="5678" heatid="25623" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="25641" lane="3" />
                <ENTRY entrytime="00:00:36.50" eventid="5694" heatid="25648" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-10-21" firstname="Lisa" gender="F" lastname="Rutkowski" nation="GER" license="377885" athleteid="23999">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.51" entrycourse="SCM" eventid="5712" heatid="25697" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.27" entrycourse="SCM" eventid="5744" heatid="25772" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:43.15" entrycourse="SCM" eventid="1123" heatid="25814" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Erem Sonsuz" gender="M" lastname="Sahin" nation="GER" license="378025" athleteid="24980">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.30" eventid="5724" heatid="25710" lane="5" />
                <ENTRY entrytime="00:01:46.57" eventid="1141" heatid="25732" lane="3" />
                <ENTRY entrytime="00:00:42.57" eventid="5740" heatid="25754" lane="2" />
                <ENTRY entrytime="00:01:45.00" eventid="7773" heatid="25781" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Jonathan" gender="M" lastname="Sandig" nation="GER" license="413757" athleteid="24220">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.34" eventid="5702" heatid="25683" lane="5" />
                <ENTRY entrytime="00:02:07.09" eventid="1141" heatid="25729" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="7773" heatid="25780" lane="6" />
                <ENTRY entrytime="00:01:41.74" eventid="1189" heatid="25829" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Diana" gender="F" lastname="Satsevich" nation="GER" license="391760" athleteid="24545">
              <ENTRIES>
                <ENTRY entrytime="00:02:55.25" eventid="1183" heatid="25672" lane="2" />
                <ENTRY entrytime="00:00:46.46" eventid="5728" heatid="25724" lane="3" />
                <ENTRY entrytime="00:01:35.90" eventid="7788" heatid="25791" lane="4" />
                <ENTRY entrytime="00:01:19.65" eventid="1195" heatid="25846" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Jan" gender="M" lastname="Schafner" nation="GER" license="406833" athleteid="24774">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1141" heatid="25730" lane="6" />
                <ENTRY entrytime="00:00:35.00" eventid="7804" heatid="25794" lane="3" />
                <ENTRY entrytime="NT" eventid="1165" heatid="25816" lane="2" />
                <ENTRY entrytime="00:02:00.00" eventid="1189" heatid="25826" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julian" gender="M" lastname="Schafner" nation="GER" license="359179" athleteid="24985">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.70" eventid="1141" heatid="25734" lane="6" />
                <ENTRY entrytime="00:00:34.92" eventid="5740" heatid="25759" lane="5" />
                <ENTRY entrytime="00:01:30.00" eventid="7773" heatid="25783" lane="2" />
                <ENTRY entrytime="00:01:19.59" eventid="1189" heatid="25833" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Maximilian" gender="M" lastname="Schechtel" nation="GER" athleteid="24779">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25607" lane="5" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25622" lane="2" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25639" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Clara" gender="F" lastname="Schiller" nation="GER" license="420943" athleteid="24550">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.24" eventid="5712" heatid="25689" lane="4" />
                <ENTRY entrytime="00:01:12.92" eventid="5728" heatid="25715" lane="2" />
                <ENTRY entrytime="00:01:02.66" eventid="5744" heatid="25762" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="7809" heatid="25798" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Elsa" gender="F" lastname="Schmaus" nation="GER" license="420936" athleteid="24555">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.15" eventid="5682" heatid="25628" lane="2" />
                <ENTRY entrytime="00:00:37.57" eventid="5698" heatid="25654" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="5664" heatid="25614" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Greta" gender="F" lastname="Schmaus" nation="GER" license="403439" athleteid="24990">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.65" eventid="5712" heatid="25695" lane="4" />
                <ENTRY entrytime="00:00:55.71" eventid="5728" heatid="25720" lane="3" />
                <ENTRY entrytime="00:01:52.52" eventid="1135" heatid="25741" lane="1" />
                <ENTRY entrytime="00:00:48.88" eventid="5744" heatid="25768" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Finja" gender="F" lastname="Schmidt" nation="GER" license="362945" athleteid="24995">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.03" eventid="5728" heatid="25725" lane="3" />
                <ENTRY entrytime="00:00:38.00" eventid="5744" heatid="25774" lane="4" />
                <ENTRY entrytime="00:01:35.00" eventid="7788" heatid="25792" lane="1" />
                <ENTRY entrytime="00:00:45.00" eventid="1123" heatid="25814" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Cem Leon" gender="M" lastname="Schulze Döring" nation="GER" license="346286" athleteid="24559">
              <ENTRIES>
                <ENTRY entrytime="00:02:39.51" eventid="1177" heatid="25664" lane="6" />
                <ENTRY entrytime="00:00:42.26" eventid="5724" heatid="25714" lane="2" />
                <ENTRY entrytime="00:01:28.09" eventid="1165" heatid="25819" lane="1" />
                <ENTRY entrytime="00:03:06.56" eventid="5655" heatid="25849" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Finn Tolgar" gender="M" lastname="Schulze Döring" nation="GER" license="368690" athleteid="24783">
              <ENTRIES>
                <ENTRY entrytime="00:01:48.00" eventid="1141" heatid="25732" lane="2" />
                <ENTRY entrytime="00:01:58.00" eventid="7773" heatid="25780" lane="1" />
                <ENTRY entrytime="00:00:48.00" eventid="1117" heatid="25807" lane="1" />
                <ENTRY entrytime="00:01:32.94" eventid="1189" heatid="25830" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Nils Ömer" gender="M" lastname="Schulze Döring" nation="GER" license="393382" athleteid="24788">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.68" eventid="1053" heatid="25611" lane="4" />
                <ENTRY entrytime="00:00:21.63" eventid="5678" heatid="25625" lane="4" />
                <ENTRY entrytime="00:00:25.03" eventid="5694" heatid="25650" lane="4" />
                <ENTRY entrytime="00:00:00.30" eventid="7701" heatid="25657" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Antonia" gender="F" lastname="Schödl" nation="GER" license="000000" athleteid="25461">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25612" lane="3" />
                <ENTRY entrytime="NT" eventid="5682" heatid="25626" lane="2" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25635" lane="1" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25651" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Julia" gender="F" lastname="Slonicz" nation="GER" license="430885" athleteid="23963">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.89" eventid="5664" heatid="25614" lane="4" />
                <ENTRY entrytime="00:00:39.55" eventid="5682" heatid="25629" lane="5" />
                <ENTRY entrytime="00:00:40.00" eventid="5690" heatid="25645" lane="1" />
                <ENTRY entrytime="00:00:39.00" eventid="5698" heatid="25654" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-11-13" firstname="Tobias" gender="M" lastname="Steger" nation="GER" athleteid="24003">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.11" entrycourse="SCM" eventid="5702" heatid="25677" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.48" entrycourse="SCM" eventid="5724" heatid="25705" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.75" entrycourse="SCM" eventid="5740" heatid="25749" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-02-19" firstname="Nick" gender="M" lastname="Steinbinder" nation="GER" athleteid="24007">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.91" entrycourse="SCM" eventid="5702" heatid="25683" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:42.86" entrycourse="SCM" eventid="5740" heatid="25754" lane="5">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25828" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Roman" gender="M" lastname="Stroh" nation="GER" license="413758" athleteid="24793">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.87" eventid="5702" heatid="25676" lane="2" />
                <ENTRY entrytime="00:01:04.16" eventid="5724" heatid="25706" lane="5" />
                <ENTRY entrytime="00:01:02.44" eventid="5740" heatid="25747" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Amir" gender="M" lastname="Tawfik" nation="GER" license="420947" athleteid="24564">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="1053" heatid="25609" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5686" heatid="25641" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Annika" gender="F" lastname="Thummerer" nation="GER" license="393378" athleteid="24225">
              <ENTRIES>
                <ENTRY entrytime="00:04:00.00" eventid="1183" heatid="25665" lane="4" />
                <ENTRY entrytime="00:02:03.40" eventid="1135" heatid="25737" lane="3" />
                <ENTRY entrytime="00:02:15.28" eventid="7788" heatid="25785" lane="2" />
                <ENTRY entrytime="00:01:56.26" eventid="1195" heatid="25838" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Carla" gender="F" lastname="Timpe" nation="GER" license="377884" athleteid="25000">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.25" eventid="5712" heatid="25695" lane="6" />
                <ENTRY entrytime="00:00:55.31" eventid="5728" heatid="25721" lane="5" />
                <ENTRY entrytime="00:00:43.61" eventid="5744" heatid="25770" lane="1" />
                <ENTRY entrytime="00:02:01.97" eventid="1135" heatid="25738" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jan" gender="M" lastname="Vilinski" nation="GER" athleteid="24567">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.00" eventid="5702" heatid="25675" lane="4" />
                <ENTRY entrytime="00:01:05.00" eventid="5724" heatid="25705" lane="3" />
                <ENTRY entrytime="00:01:02.00" eventid="5740" heatid="25748" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-04" firstname="Emily" gender="F" lastname="Wech" nation="GER" license="359178" athleteid="24011">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.07" entrycourse="SCM" eventid="1135" heatid="25741" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.74" entrycourse="SCM" eventid="7788" heatid="25788" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.71" entrycourse="SCM" eventid="1171" heatid="25820" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leander" gender="M" lastname="Wech" nation="GER" license="392571" athleteid="24571">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.85" eventid="5702" heatid="25675" lane="1" />
                <ENTRY entrytime="00:01:08.33" eventid="5724" heatid="25705" lane="6" />
                <ENTRY entrytime="00:01:02.39" eventid="5740" heatid="25747" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="7804" heatid="25794" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-10-19" firstname="Patrick" gender="M" lastname="Wech" nation="GER" license="392572" athleteid="24015">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.08" entrycourse="SCM" eventid="5724" heatid="25710" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-11-10" name="42. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.05" entrycourse="SCM" eventid="5740" heatid="25753" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.77" entrycourse="SCM" eventid="1117" heatid="25805" lane="1">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Anna-Lena" gender="F" lastname="Weisbrodt" nation="GER" license="407277" athleteid="25005">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.00" eventid="5712" heatid="25695" lane="3" />
                <ENTRY entrytime="00:00:45.00" eventid="5728" heatid="25726" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5744" heatid="25766" lane="3" />
                <ENTRY entrytime="00:01:55.00" eventid="1171" heatid="25821" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Benjamin" gender="M" lastname="Welker" nation="GER" license="392569" athleteid="23968">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.56" eventid="5724" heatid="25707" lane="4" />
                <ENTRY entrytime="00:02:15.00" eventid="1141" heatid="25729" lane="5" />
                <ENTRY entrytime="00:00:25.00" eventid="7804" heatid="25797" lane="5" />
                <ENTRY entrytime="00:02:15.00" eventid="1189" heatid="25825" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Henri" gender="M" lastname="Wittl" nation="GER" athleteid="23973">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1053" heatid="25608" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="7691" heatid="25632" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25640" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julia" gender="F" lastname="Wolf" nation="GER" license="362947" athleteid="24576">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.15" eventid="1111" heatid="25703" lane="4" />
                <ENTRY entrytime="00:01:44.43" eventid="1135" heatid="25743" lane="3" />
                <ENTRY entrytime="00:01:32.82" eventid="7788" heatid="25792" lane="3" />
                <ENTRY entrytime="00:01:18.97" eventid="1195" heatid="25847" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Jan" gender="M" lastname="Zeidler" nation="GER" license="389378" athleteid="24797">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5702" heatid="25677" lane="3" />
                <ENTRY entrytime="NT" eventid="5724" heatid="25704" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="25749" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2015-01-01" firstname="Simon" gender="M" lastname="Zeidler" nation="GER" license="0" athleteid="24801">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.27" eventid="1053" heatid="25608" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="5678" heatid="25622" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25640" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-04-24" firstname="Arijalda" gender="F" lastname="Zukorlic" nation="GER" athleteid="24019">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25685" lane="2" />
                <ENTRY entrytime="NT" eventid="5728" heatid="25715" lane="6" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25761" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5085" nation="GER" region="02" clubid="24333" name="SG Bamberg">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="Elias" gender="M" lastname="Becker" nation="GER" license="429038" athleteid="24334">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="5702" heatid="25673" lane="4" />
                <ENTRY entrytime="00:01:20.00" eventid="5740" heatid="25747" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Katharina" gender="F" lastname="Dieter" nation="GER" license="0" athleteid="24337">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="25626" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25636" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="25644" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Sanja" gender="F" lastname="Dietzel" nation="GER" license="0" athleteid="24341">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="25628" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25636" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Mara" gender="F" lastname="Friedemann" nation="GER" license="434413" athleteid="24344">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.00" eventid="5712" heatid="25686" lane="5" />
                <ENTRY entrytime="00:01:30.00" eventid="5744" heatid="25761" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Leo" gender="M" lastname="Gebhard" nation="GER" license="425301" athleteid="24347">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.11" eventid="5702" heatid="25674" lane="6" />
                <ENTRY entrytime="00:01:10.00" eventid="5724" heatid="25704" lane="3" />
                <ENTRY entrytime="00:00:58.76" eventid="5740" heatid="25749" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Elisa" gender="F" lastname="Graf" nation="GER" license="0" athleteid="24351">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.94" eventid="5664" heatid="25613" lane="3" />
                <ENTRY entrytime="00:00:43.73" eventid="5682" heatid="25629" lane="6" />
                <ENTRY entrytime="00:00:55.00" eventid="7696" heatid="25636" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Emilia" gender="F" lastname="Graf" nation="GER" license="429036" athleteid="24355">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.00" eventid="5712" heatid="25686" lane="3" />
                <ENTRY entrytime="00:01:12.00" eventid="5728" heatid="25715" lane="4" />
                <ENTRY entrytime="00:01:06.00" eventid="5744" heatid="25762" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Moritz" gender="M" lastname="Hartmann" nation="GER" license="0" athleteid="24359">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.00" eventid="1053" heatid="25608" lane="2" />
                <ENTRY entrytime="00:00:50.00" eventid="5678" heatid="25623" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="7691" heatid="25632" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25639" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Juna" gender="F" lastname="Heinze" nation="GER" license="0" athleteid="24364">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="25627" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Paula" gender="F" lastname="Heinze" nation="GER" license="395455" athleteid="24366">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.00" eventid="5712" heatid="25687" lane="3" />
                <ENTRY entrytime="00:01:09.00" eventid="5728" heatid="25716" lane="1" />
                <ENTRY entrytime="00:00:59.10" eventid="5744" heatid="25764" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Jannik" gender="M" lastname="Hünniger" nation="GER" license="409224" athleteid="24370">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.78" eventid="5702" heatid="25682" lane="1" />
                <ENTRY entrytime="00:00:47.54" eventid="5724" heatid="25712" lane="4" />
                <ENTRY entrytime="00:01:41.37" eventid="7773" heatid="25781" lane="3" />
                <ENTRY entrytime="00:01:46.00" eventid="1165" heatid="25817" lane="1" />
                <ENTRY entrytime="00:01:30.99" eventid="1189" heatid="25831" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lara" gender="F" lastname="Hünniger" nation="GER" license="425312" athleteid="24376">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.00" eventid="5712" heatid="25687" lane="6" />
                <ENTRY entrytime="00:00:59.20" eventid="5744" heatid="25763" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Timurs" gender="M" lastname="Iljins" nation="GER" license="409220" athleteid="24379">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="5702" heatid="25673" lane="3" />
                <ENTRY entrytime="00:00:58.88" eventid="5724" heatid="25707" lane="2" />
                <ENTRY entrytime="00:00:48.93" eventid="5740" heatid="25751" lane="3" />
                <ENTRY entrytime="00:02:15.00" eventid="7773" heatid="25778" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Eva" gender="F" lastname="Jakubaß" nation="GER" license="409223" athleteid="24384">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.80" eventid="5712" heatid="25688" lane="3" />
                <ENTRY entrytime="00:00:55.18" eventid="5728" heatid="25721" lane="2" />
                <ENTRY entrytime="00:00:48.65" eventid="5744" heatid="25768" lane="5" />
                <ENTRY entrytime="00:01:48.08" eventid="1195" heatid="25840" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Raphael" gender="M" lastname="Jakubaß" nation="GER" license="392827" athleteid="24389">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.99" eventid="5702" heatid="25678" lane="3" />
                <ENTRY entrytime="00:00:43.27" eventid="5740" heatid="25754" lane="1" />
                <ENTRY entrytime="00:01:50.00" eventid="7773" heatid="25780" lane="4" />
                <ENTRY entrytime="00:00:48.70" eventid="1117" heatid="25806" lane="3" />
                <ENTRY entrytime="00:01:39.77" eventid="1189" heatid="25829" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Sebastian" gender="M" lastname="Jakubaß" nation="GER" license="0" athleteid="24395">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5678" heatid="25623" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="7691" heatid="25633" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25640" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Antonio" gender="M" lastname="La Corte" nation="GER" license="0" athleteid="24399">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5678" heatid="25623" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25640" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Olivia" gender="F" lastname="Lang" nation="GER" license="425304" athleteid="24402">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5728" heatid="25715" lane="3" />
                <ENTRY entrytime="00:01:01.82" eventid="5744" heatid="25763" lane="6" />
                <ENTRY entrytime="00:00:36.00" eventid="7809" heatid="25798" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Samuel" gender="M" lastname="Lang" nation="GER" license="392828" athleteid="24406">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.00" eventid="1177" heatid="25662" lane="1" />
                <ENTRY entrytime="00:01:46.84" eventid="1103" heatid="25699" lane="5" />
                <ENTRY entrytime="00:00:37.28" eventid="5740" heatid="25758" lane="6" />
                <ENTRY entrytime="00:00:44.10" eventid="1117" heatid="25807" lane="4" />
                <ENTRY entrytime="00:01:25.60" eventid="1189" heatid="25833" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Eva" gender="F" lastname="Meister" nation="GER" license="409222" athleteid="24412">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.62" eventid="5712" heatid="25694" lane="6" />
                <ENTRY entrytime="00:01:02.76" eventid="5728" heatid="25717" lane="1" />
                <ENTRY entrytime="00:00:48.90" eventid="5744" heatid="25767" lane="3" />
                <ENTRY entrytime="00:02:07.00" eventid="7788" heatid="25786" lane="1" />
                <ENTRY entrytime="00:00:32.00" eventid="7809" heatid="25799" lane="5" />
                <ENTRY entrytime="00:01:55.00" eventid="1195" heatid="25838" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Jakob" gender="M" lastname="Meister" nation="GER" license="361866" athleteid="24419">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.00" eventid="5702" heatid="25683" lane="1" />
                <ENTRY entrytime="00:00:45.00" eventid="5724" heatid="25713" lane="3" />
                <ENTRY entrytime="00:00:38.00" eventid="5740" heatid="25757" lane="4" />
                <ENTRY entrytime="00:00:47.00" eventid="1117" heatid="25807" lane="5" />
                <ENTRY entrytime="00:01:39.00" eventid="1165" heatid="25818" lane="6" />
                <ENTRY entrytime="00:03:30.00" eventid="5655" heatid="25848" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Paul" gender="M" lastname="Nitsche" nation="GER" license="434412" athleteid="24426">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.00" eventid="5702" heatid="25673" lane="1" />
                <ENTRY entrytime="00:01:30.00" eventid="5740" heatid="25746" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Noa-Louis" gender="M" lastname="Panknin" nation="GER" license="429039" athleteid="24429">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5702" heatid="25674" lane="5" />
                <ENTRY entrytime="00:01:10.00" eventid="5740" heatid="25747" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Linda" gender="F" lastname="Schellenberger" nation="GER" license="0" athleteid="24432">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.00" eventid="5674" heatid="25621" lane="3" />
                <ENTRY entrytime="00:00:24.92" eventid="5682" heatid="25631" lane="4" />
                <ENTRY entrytime="00:00:29.10" eventid="7696" heatid="25638" lane="3" />
                <ENTRY entrytime="00:00:28.25" eventid="5698" heatid="25656" lane="2" />
                <ENTRY entrytime="00:00:36.00" eventid="7706" heatid="25658" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Marie" gender="F" lastname="Schellenberger" nation="GER" license="0" athleteid="24438">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.40" eventid="5664" heatid="25616" lane="4" />
                <ENTRY entrytime="00:00:33.06" eventid="5682" heatid="25630" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" heatid="25637" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5690" heatid="25644" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lara" gender="F" lastname="Schindler" nation="GER" license="409221" athleteid="24443">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.26" eventid="5712" heatid="25692" lane="3" />
                <ENTRY entrytime="00:00:59.28" eventid="5728" heatid="25720" lane="1" />
                <ENTRY entrytime="00:00:52.03" eventid="5744" heatid="25765" lane="3" />
                <ENTRY entrytime="00:02:07.00" eventid="7788" heatid="25786" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Luisa" gender="F" lastname="Schindler" nation="GER" license="0" athleteid="24448">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5664" heatid="25613" lane="5" />
                <ENTRY entrytime="00:00:57.46" eventid="5682" heatid="25628" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25635" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Paula" gender="F" lastname="Schuh" nation="GER" license="425299" athleteid="24452">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.11" eventid="5712" heatid="25689" lane="5" />
                <ENTRY entrytime="00:01:09.00" eventid="5728" heatid="25716" lane="5" />
                <ENTRY entrytime="00:00:56.49" eventid="5744" heatid="25764" lane="1" />
                <ENTRY entrytime="00:02:10.00" eventid="7788" heatid="25785" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Hanna" gender="F" lastname="Skamrahl" nation="GER" license="0" athleteid="24457">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5664" heatid="25613" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="25627" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="25643" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Antonia" gender="F" lastname="Struckmeier" nation="GER" license="0" athleteid="24461">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.36" eventid="5664" heatid="25614" lane="1" />
                <ENTRY entrytime="00:00:44.00" eventid="5674" heatid="25621" lane="4" />
                <ENTRY entrytime="00:00:32.20" eventid="5682" heatid="25630" lane="2" />
                <ENTRY entrytime="00:00:36.90" eventid="7696" heatid="25638" lane="2" />
                <ENTRY entrytime="00:00:41.34" eventid="5698" heatid="25654" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Troll" nation="GER" license="0" athleteid="24467">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5664" heatid="25613" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="25627" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25636" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lilia" gender="F" lastname="Wagner" nation="GER" license="0" athleteid="24471">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="25627" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25635" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="25644" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Laurin" gender="M" lastname="Willenberg" nation="GER" license="430362" athleteid="24475">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="5702" heatid="25673" lane="2" />
                <ENTRY entrytime="00:01:20.00" eventid="5740" heatid="25747" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Fiona" gender="F" lastname="Wystrach" nation="GER" license="0" athleteid="24478">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5682" heatid="25627" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25636" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="25644" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="5095" nation="GER" region="02" clubid="24581" name="SG Frankenhöhe">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="Laura" gender="F" lastname="Bauereiß" nation="GER" license="000000" athleteid="24582">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.00" eventid="5712" heatid="25692" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25718" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5744" heatid="25766" lane="2" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25798" lane="6" />
                <ENTRY entrytime="00:02:10.00" eventid="1195" heatid="25836" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Noah" gender="M" lastname="Binder" nation="GER" license="000000" athleteid="24588">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.00" eventid="5702" heatid="25681" lane="3" />
                <ENTRY entrytime="00:00:54.00" eventid="5724" heatid="25709" lane="4" />
                <ENTRY entrytime="00:00:39.00" eventid="5740" heatid="25756" lane="4" />
                <ENTRY entrytime="00:00:55.00" eventid="1117" heatid="25805" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Antonia" gender="F" lastname="Bößendorfer" nation="GER" license="364988" athleteid="24593">
              <ENTRIES>
                <ENTRY entrytime="00:03:01.27" eventid="1183" heatid="25671" lane="4" />
                <ENTRY entrytime="00:01:50.00" eventid="1135" heatid="25742" lane="6" />
                <ENTRY entrytime="00:00:37.00" eventid="5744" heatid="25775" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="1123" heatid="25812" lane="1" />
                <ENTRY entrytime="00:01:25.00" eventid="1195" heatid="25845" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Emely" gender="F" lastname="Bößendörfer" nation="GER" license="364989" athleteid="24599">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.00" eventid="1183" heatid="25671" lane="5" />
                <ENTRY entrytime="00:01:40.00" eventid="1135" heatid="25744" lane="2" />
                <ENTRY entrytime="00:00:36.00" eventid="5744" heatid="25776" lane="1" />
                <ENTRY entrytime="00:00:44.00" eventid="1123" heatid="25814" lane="4" />
                <ENTRY entrytime="00:01:23.00" eventid="1195" heatid="25845" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Anne" gender="F" lastname="Frank" nation="GER" license="000000" athleteid="24605">
              <ENTRIES>
                <ENTRY entrytime="00:03:22.00" eventid="1183" heatid="25669" lane="4" />
                <ENTRY entrytime="00:01:49.00" eventid="1135" heatid="25742" lane="4" />
                <ENTRY entrytime="00:00:39.00" eventid="5744" heatid="25773" lane="4" />
                <ENTRY entrytime="00:00:55.00" eventid="1123" heatid="25810" lane="4" />
                <ENTRY entrytime="00:01:34.00" eventid="1195" heatid="25842" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lana" gender="F" lastname="Freisler" nation="GER" license="392397" athleteid="24611">
              <ENTRIES>
                <ENTRY entrytime="00:03:14.00" eventid="1183" heatid="25670" lane="3" />
                <ENTRY entrytime="00:01:45.00" eventid="1135" heatid="25743" lane="4" />
                <ENTRY entrytime="00:00:41.00" eventid="5744" heatid="25771" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="1123" heatid="25812" lane="6" />
                <ENTRY entrytime="00:01:32.00" eventid="1195" heatid="25842" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Jonah" gender="M" lastname="Henninger" nation="GER" license="379527" athleteid="24617">
              <ENTRIES>
                <ENTRY entrytime="00:02:25.00" eventid="1177" heatid="25664" lane="2" />
                <ENTRY entrytime="00:01:20.00" eventid="1103" heatid="25700" lane="3" />
                <ENTRY entrytime="00:00:29.00" eventid="5740" heatid="25760" lane="3" />
                <ENTRY entrytime="00:01:24.00" eventid="1165" heatid="25819" lane="5" />
                <ENTRY entrytime="00:01:05.00" eventid="1189" heatid="25835" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lea" gender="F" lastname="Herrmann" nation="GER" license="000000" athleteid="24623">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.00" eventid="5712" heatid="25693" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25718" lane="1" />
                <ENTRY entrytime="00:00:49.00" eventid="5744" heatid="25767" lane="5" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25798" lane="1" />
                <ENTRY entrytime="00:01:55.00" eventid="1195" heatid="25838" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Hanna" gender="F" lastname="Kachelrieß" nation="GER" license="392395" athleteid="24629">
              <ENTRIES>
                <ENTRY entrytime="00:03:25.00" eventid="1183" heatid="25669" lane="6" />
                <ENTRY entrytime="00:01:51.00" eventid="1135" heatid="25741" lane="3" />
                <ENTRY entrytime="00:00:39.00" eventid="5744" heatid="25773" lane="3" />
                <ENTRY entrytime="00:00:55.00" eventid="1123" heatid="25810" lane="3" />
                <ENTRY entrytime="00:01:31.00" eventid="1195" heatid="25843" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Julia" gender="F" lastname="KLaußecker" nation="GER" license="000000" athleteid="24635">
              <ENTRIES>
                <ENTRY entrytime="00:04:00.00" eventid="1183" heatid="25665" lane="3" />
                <ENTRY entrytime="00:01:55.00" eventid="1135" heatid="25740" lane="4" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="25765" lane="6" />
                <ENTRY entrytime="00:02:05.00" eventid="1195" heatid="25837" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Sophia" gender="F" lastname="Kloha" nation="GER" license="000000" athleteid="24639">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.00" eventid="5712" heatid="25691" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25718" lane="2" />
                <ENTRY entrytime="00:00:49.00" eventid="5744" heatid="25767" lane="4" />
                <ENTRY entrytime="00:01:55.00" eventid="1195" heatid="25838" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Eleni" gender="F" lastname="Martin" nation="GER" license="000000" athleteid="24644">
              <ENTRIES>
                <ENTRY entrytime="00:03:35.00" eventid="1183" heatid="25667" lane="3" />
                <ENTRY entrytime="00:01:55.00" eventid="1135" heatid="25740" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="5744" heatid="25772" lane="4" />
                <ENTRY entrytime="00:01:38.00" eventid="1195" heatid="25841" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Eileen" gender="F" lastname="Möhring" nation="GER" license="000000" athleteid="24649">
              <ENTRIES>
                <ENTRY entrytime="00:02:58.00" eventid="1183" heatid="25672" lane="6" />
                <ENTRY entrytime="00:00:48.00" eventid="5728" heatid="25724" lane="6" />
                <ENTRY entrytime="00:00:36.00" eventid="5744" heatid="25776" lane="5" />
                <ENTRY entrytime="00:01:25.00" eventid="1195" heatid="25845" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Tilly" gender="F" lastname="Neumeyer" nation="GER" license="000000" athleteid="24654">
              <ENTRIES>
                <ENTRY entrytime="00:03:50.00" eventid="1183" heatid="25666" lane="4" />
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="25738" lane="2" />
                <ENTRY entrytime="00:00:45.00" eventid="5744" heatid="25769" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="1195" heatid="25839" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Laurens" gender="M" lastname="Springer" nation="GER" license="000000" athleteid="24659">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.00" eventid="5702" heatid="25675" lane="3" />
                <ENTRY entrytime="00:01:08.00" eventid="5724" heatid="25705" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="5740" heatid="25751" lane="6" />
                <ENTRY entrytime="00:01:55.00" eventid="1189" heatid="25827" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6768" nation="GER" region="02" clubid="25010" name="SG Mittelfranken">
          <ATHLETES>
            <ATHLETE birthdate="2006-01-01" firstname="Paulina" gender="F" lastname="Artavia" nation="GER" license="377714" athleteid="25011">
              <ENTRIES>
                <ENTRY entrytime="00:03:20.19" eventid="1183" heatid="25669" lane="3" />
                <ENTRY entrytime="00:00:38.74" eventid="5728" heatid="25727" lane="4" />
                <ENTRY entrytime="00:01:39.75" eventid="1135" heatid="25744" lane="3" />
                <ENTRY entrytime="00:01:29.59" eventid="7788" heatid="25793" lane="2" />
                <ENTRY entrytime="00:01:24.18" eventid="1171" heatid="25824" lane="4" />
                <ENTRY entrytime="00:01:22.78" eventid="1195" heatid="25846" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Liv" gender="F" lastname="Asse" nation="GER" license="406748" athleteid="25018">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.95" eventid="5712" heatid="25696" lane="6" />
                <ENTRY entrytime="00:01:55.62" eventid="1135" heatid="25740" lane="1" />
                <ENTRY entrytime="00:01:53.01" eventid="7788" heatid="25788" lane="4" />
                <ENTRY entrytime="00:00:47.62" eventid="1123" heatid="25813" lane="5" />
                <ENTRY entrytime="00:01:46.47" eventid="1171" heatid="25822" lane="6" />
                <ENTRY entrytime="00:01:31.71" eventid="1195" heatid="25843" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emelie" gender="F" lastname="Bachmeier" nation="GER" license="432643" athleteid="25025">
              <ENTRIES>
                <ENTRY entrytime="00:03:15.00" eventid="1183" heatid="25670" lane="4" />
                <ENTRY entrytime="00:00:41.00" eventid="5728" heatid="25727" lane="1" />
                <ENTRY entrytime="00:00:38.50" eventid="5744" heatid="25774" lane="1" />
                <ENTRY entrytime="00:01:35.00" eventid="7788" heatid="25792" lane="6" />
                <ENTRY entrytime="00:00:48.00" eventid="1123" heatid="25812" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Alexandra" gender="F" lastname="Banosopoulou" nation="GER" license="417319" athleteid="25031">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.16" eventid="5664" heatid="25617" lane="2" />
                <ENTRY entrytime="00:00:23.97" eventid="5682" heatid="25631" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="7696" heatid="25638" lane="4" />
                <ENTRY entrytime="00:00:35.00" eventid="5690" heatid="25646" lane="1" />
                <ENTRY entrytime="00:00:26.90" eventid="5698" heatid="25656" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Freyja" gender="F" lastname="Bay" nation="GER" license="0" athleteid="25037">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.00" eventid="5664" heatid="25617" lane="3" />
                <ENTRY entrytime="00:00:25.00" eventid="5682" heatid="25631" lane="5" />
                <ENTRY entrytime="00:00:32.00" eventid="5690" heatid="25646" lane="2" />
                <ENTRY entrytime="00:00:25.00" eventid="5698" heatid="25656" lane="3" />
                <ENTRY entrytime="00:00:40.00" eventid="7706" heatid="25658" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Stella" gender="F" lastname="Bay" nation="GER" license="427351" athleteid="25043">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.00" eventid="5712" heatid="25693" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25719" lane="6" />
                <ENTRY entrytime="00:00:54.00" eventid="5744" heatid="25765" lane="4" />
                <ENTRY entrytime="00:00:28.50" eventid="7809" heatid="25800" lane="4" />
                <ENTRY entrytime="00:02:08.00" eventid="1195" heatid="25837" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Sebastian" gender="M" lastname="Brandner" nation="GER" license="406001" athleteid="25049">
              <ENTRIES>
                <ENTRY entrytime="00:03:39.14" eventid="1177" heatid="25660" lane="5" />
                <ENTRY entrytime="00:00:54.62" eventid="5702" heatid="25680" lane="1" />
                <ENTRY entrytime="00:01:37.11" eventid="7773" heatid="25782" lane="2" />
                <ENTRY entrytime="00:00:49.09" eventid="1117" heatid="25806" lane="4" />
                <ENTRY entrytime="00:01:26.40" eventid="1189" heatid="25832" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Pia" gender="F" lastname="Braun" nation="GER" license="383927" athleteid="25055">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.43" eventid="5712" heatid="25698" lane="5" />
                <ENTRY entrytime="00:00:44.78" eventid="5728" heatid="25726" lane="1" />
                <ENTRY entrytime="00:01:40.40" eventid="1135" heatid="25744" lane="5" />
                <ENTRY entrytime="00:01:37.50" eventid="7788" heatid="25791" lane="2" />
                <ENTRY entrytime="00:01:40.53" eventid="1171" heatid="25823" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Isabelle Zoe" gender="F" lastname="Brauns" nation="GER" license="415616" athleteid="25061">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.02" eventid="5712" heatid="25694" lane="4" />
                <ENTRY entrytime="00:00:46.59" eventid="5728" heatid="25724" lane="4" />
                <ENTRY entrytime="00:00:45.60" eventid="5744" heatid="25769" lane="5" />
                <ENTRY entrytime="00:00:49.16" eventid="1123" heatid="25812" lane="5" />
                <ENTRY entrytime="00:03:45.00" eventid="5661" heatid="25850" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Helena" gender="F" lastname="Brausam" nation="GER" license="420240" athleteid="25067">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.59" eventid="5712" heatid="25694" lane="3" />
                <ENTRY entrytime="00:02:10.09" eventid="1135" heatid="25736" lane="4" />
                <ENTRY entrytime="00:00:59.75" eventid="5744" heatid="25763" lane="4" />
                <ENTRY entrytime="00:02:00.00" eventid="1195" heatid="25838" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Marie" gender="F" lastname="Brunner" nation="GER" license="417323" athleteid="25072">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.31" eventid="5712" heatid="25690" lane="1" />
                <ENTRY entrytime="00:00:55.59" eventid="5728" heatid="25721" lane="1" />
                <ENTRY entrytime="00:00:47.94" eventid="5744" heatid="25768" lane="2" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25801" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Emilia" gender="F" lastname="Burdack" nation="GER" license="417324" athleteid="25077">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.47" eventid="5712" heatid="25694" lane="1" />
                <ENTRY entrytime="00:01:00.96" eventid="5728" heatid="25718" lane="6" />
                <ENTRY entrytime="00:00:49.72" eventid="5744" heatid="25767" lane="6" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25802" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Paul Wilfried Jens" gender="M" lastname="Burkhardt" nation="GER" license="406751" athleteid="25082">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.90" eventid="5702" heatid="25674" lane="3" />
                <ENTRY entrytime="00:00:50.84" eventid="5724" heatid="25710" lane="4" />
                <ENTRY entrytime="00:00:55.45" eventid="5740" heatid="25750" lane="1" />
                <ENTRY entrytime="00:02:00.00" eventid="7773" heatid="25779" lane="3" />
                <ENTRY entrytime="00:01:54.16" eventid="1165" heatid="25816" lane="3" />
                <ENTRY entrytime="00:01:50.47" eventid="1189" heatid="25827" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Anton" gender="M" lastname="Cao" nation="GER" license="417199" athleteid="25089">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.12" eventid="5702" heatid="25681" lane="1" />
                <ENTRY entrytime="00:00:51.35" eventid="5724" heatid="25710" lane="2" />
                <ENTRY entrytime="00:00:42.30" eventid="5740" heatid="25754" lane="4" />
                <ENTRY entrytime="00:00:25.00" eventid="7804" heatid="25796" lane="4" />
                <ENTRY entrytime="00:01:46.46" eventid="1189" heatid="25828" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Kai" gender="M" lastname="Chan" nation="GER" license="392890" athleteid="25095">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.24" eventid="5702" heatid="25681" lane="4" />
                <ENTRY entrytime="00:00:48.13" eventid="5724" heatid="25712" lane="1" />
                <ENTRY entrytime="00:01:50.99" eventid="1141" heatid="25731" lane="3" />
                <ENTRY entrytime="00:00:40.53" eventid="5740" heatid="25756" lane="6" />
                <ENTRY entrytime="00:01:43.34" eventid="1165" heatid="25817" lane="2" />
                <ENTRY entrytime="00:01:35.56" eventid="1189" heatid="25830" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Stefan" gender="M" lastname="David" nation="GER" license="0" athleteid="25102">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.00" eventid="1053" heatid="25611" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="5668" heatid="25619" lane="4" />
                <ENTRY entrytime="00:00:25.00" eventid="5678" heatid="25625" lane="2" />
                <ENTRY entrytime="00:00:35.00" eventid="7691" heatid="25634" lane="2" />
                <ENTRY entrytime="00:00:25.00" eventid="5694" heatid="25650" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Timur" gender="M" lastname="Dick" nation="GER" license="420056" athleteid="25108">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.65" eventid="5702" heatid="25675" lane="5" />
                <ENTRY entrytime="00:01:02.34" eventid="5724" heatid="25706" lane="2" />
                <ENTRY entrytime="00:00:57.66" eventid="5740" heatid="25749" lane="3" />
                <ENTRY entrytime="00:00:25.00" eventid="7804" heatid="25797" lane="6" />
                <ENTRY entrytime="00:02:08.00" eventid="1189" heatid="25826" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="David" gender="M" lastname="Engler" nation="GER" license="406755" athleteid="25114">
              <ENTRIES>
                <ENTRY entrytime="00:03:18.08" eventid="1177" heatid="25661" lane="5" />
                <ENTRY entrytime="00:00:45.69" eventid="5702" heatid="25683" lane="2" />
                <ENTRY entrytime="00:01:35.34" eventid="1141" heatid="25733" lane="3" />
                <ENTRY entrytime="00:00:49.36" eventid="1117" heatid="25806" lane="2" />
                <ENTRY entrytime="00:01:38.77" eventid="1165" heatid="25818" lane="1" />
                <ENTRY entrytime="00:01:27.12" eventid="1189" heatid="25832" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Daniel" gender="M" lastname="Frank" nation="GER" license="0" athleteid="25121">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="1053" heatid="25609" lane="1" />
                <ENTRY entrytime="00:00:40.00" eventid="5678" heatid="25623" lane="2" />
                <ENTRY entrytime="00:00:45.00" eventid="7691" heatid="25633" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="5686" heatid="25641" lane="5" />
                <ENTRY entrytime="00:00:40.00" eventid="5694" heatid="25648" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Peter" gender="M" lastname="Grießinger" nation="GER" license="377882" athleteid="25348">
              <ENTRIES>
                <ENTRY entrytime="00:03:15.00" eventid="1177" heatid="25661" lane="3" />
                <ENTRY entrytime="00:01:55.00" eventid="1141" heatid="25731" lane="4" />
                <ENTRY entrytime="00:01:50.00" eventid="7773" heatid="25781" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="1117" heatid="25805" lane="6" />
                <ENTRY entrytime="00:01:40.00" eventid="1165" heatid="25817" lane="3" />
                <ENTRY entrytime="00:01:30.00" eventid="1189" heatid="25831" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Arthur" gender="M" lastname="Gross" nation="GER" license="420054" athleteid="25127">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.60" eventid="5702" heatid="25676" lane="6" />
                <ENTRY entrytime="00:00:49.15" eventid="5724" heatid="25711" lane="4" />
                <ENTRY entrytime="00:00:40.80" eventid="5740" heatid="25755" lane="4" />
                <ENTRY entrytime="00:00:51.60" eventid="1117" heatid="25806" lane="6" />
                <ENTRY entrytime="00:01:36.12" eventid="1189" heatid="25830" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Roman" gender="M" lastname="Gross" nation="GER" license="420055" athleteid="25133">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.82" eventid="5702" heatid="25677" lane="1" />
                <ENTRY entrytime="00:00:48.22" eventid="5724" heatid="25712" lane="6" />
                <ENTRY entrytime="00:00:38.54" eventid="5740" heatid="25757" lane="6" />
                <ENTRY entrytime="00:00:49.36" eventid="1117" heatid="25806" lane="5" />
                <ENTRY entrytime="00:03:35.00" eventid="5655" heatid="25848" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Julian" gender="M" lastname="Hampel" nation="GER" license="401463" athleteid="25139">
              <ENTRIES>
                <ENTRY entrytime="00:03:22.06" eventid="1177" heatid="25661" lane="1" />
                <ENTRY entrytime="00:00:43.61" eventid="5724" heatid="25714" lane="5" />
                <ENTRY entrytime="00:01:52.68" eventid="7773" heatid="25780" lane="2" />
                <ENTRY entrytime="00:00:42.23" eventid="1117" heatid="25808" lane="1" />
                <ENTRY entrytime="00:01:24.45" eventid="1189" heatid="25833" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Helena" gender="F" lastname="Hauer" nation="GER" license="406750" athleteid="25145">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.96" eventid="5712" heatid="25693" lane="3" />
                <ENTRY entrytime="00:00:45.91" eventid="5728" heatid="25725" lane="2" />
                <ENTRY entrytime="00:00:40.44" eventid="5744" heatid="25771" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="1123" heatid="25809" lane="2" />
                <ENTRY entrytime="00:01:41.06" eventid="1171" heatid="25822" lane="4" />
                <ENTRY entrytime="00:01:34.32" eventid="1195" heatid="25841" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Eymen" gender="M" lastname="Hayirli" nation="GER" license="414887" athleteid="25152">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.10" eventid="1053" heatid="25611" lane="1" />
                <ENTRY entrytime="00:00:30.00" eventid="5668" heatid="25619" lane="3" />
                <ENTRY entrytime="00:00:20.20" eventid="5678" heatid="25625" lane="3" />
                <ENTRY entrytime="00:00:30.00" eventid="5686" heatid="25642" lane="5" />
                <ENTRY entrytime="00:00:27.75" eventid="5694" heatid="25650" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Hanna" gender="F" lastname="Holtmannspötter" nation="GER" license="420811" athleteid="25158">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.31" eventid="5712" heatid="25686" lane="2" />
                <ENTRY entrytime="00:01:06.05" eventid="5728" heatid="25716" lane="4" />
                <ENTRY entrytime="00:00:47.56" eventid="5744" heatid="25768" lane="4" />
                <ENTRY entrytime="00:02:10.00" eventid="1195" heatid="25836" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lilly" gender="F" lastname="Jeschke" nation="GER" license="427348" athleteid="25163">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5712" heatid="25690" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25719" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25763" lane="5" />
                <ENTRY entrytime="00:00:30.00" eventid="7809" heatid="25800" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Anna-Lena" gender="F" lastname="Karasek" nation="GER" license="418668" athleteid="25168">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.03" eventid="5664" heatid="25617" lane="5" />
                <ENTRY entrytime="00:00:29.67" eventid="5682" heatid="25631" lane="6" />
                <ENTRY entrytime="00:00:30.00" eventid="5690" heatid="25646" lane="4" />
                <ENTRY entrytime="00:00:28.72" eventid="5698" heatid="25656" lane="5" />
                <ENTRY entrytime="00:00:35.00" eventid="7706" heatid="25658" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Laura" gender="F" lastname="Kim" nation="GER" license="417320" athleteid="25174">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.34" eventid="5712" heatid="25688" lane="5" />
                <ENTRY entrytime="00:00:59.81" eventid="5728" heatid="25719" lane="3" />
                <ENTRY entrytime="00:00:55.82" eventid="5744" heatid="25764" lane="5" />
                <ENTRY entrytime="00:00:30.00" eventid="7809" heatid="25799" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Ella" gender="F" lastname="Kleinert" nation="GER" license="412139" athleteid="25179">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.51" eventid="5712" heatid="25692" lane="2" />
                <ENTRY entrytime="00:00:53.31" eventid="5728" heatid="25722" lane="6" />
                <ENTRY entrytime="00:00:49.33" eventid="5744" heatid="25767" lane="1" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25801" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="1195" heatid="25839" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jonathan" gender="M" lastname="Koepnick" nation="GER" license="408297" athleteid="25185">
              <ENTRIES>
                <ENTRY entrytime="00:01:44.26" eventid="1103" heatid="25699" lane="4" />
                <ENTRY entrytime="00:00:35.86" eventid="5740" heatid="25758" lane="4" />
                <ENTRY entrytime="00:01:27.30" eventid="7773" heatid="25784" lane="1" />
                <ENTRY entrytime="00:00:43.53" eventid="1117" heatid="25808" lane="6" />
                <ENTRY entrytime="00:01:28.32" eventid="1165" heatid="25819" lane="6" />
                <ENTRY entrytime="00:01:17.53" eventid="1189" heatid="25834" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Dennis" gender="M" lastname="Kranz" nation="GER" license="425761" athleteid="25231">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="1053" heatid="25609" lane="3" />
                <ENTRY entrytime="00:00:31.00" eventid="5678" heatid="25624" lane="4" />
                <ENTRY entrytime="00:00:40.00" eventid="7691" heatid="25634" lane="6" />
                <ENTRY entrytime="00:00:35.00" eventid="5686" heatid="25642" lane="6" />
                <ENTRY entrytime="00:00:40.00" eventid="5694" heatid="25647" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Alessia" gender="F" lastname="Köhler" nation="GER" license="399200" athleteid="25192">
              <ENTRIES>
                <ENTRY entrytime="00:02:55.98" eventid="1183" heatid="25672" lane="5" />
                <ENTRY entrytime="00:01:36.05" eventid="1111" heatid="25703" lane="2" />
                <ENTRY entrytime="00:00:44.70" eventid="5728" heatid="25726" lane="2" />
                <ENTRY entrytime="00:01:33.60" eventid="7788" heatid="25792" lane="4" />
                <ENTRY entrytime="00:01:21.31" eventid="1195" heatid="25846" lane="1" />
                <ENTRY entrytime="00:03:15.43" eventid="5661" heatid="25851" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ida" gender="F" lastname="Köhler" nation="GER" license="428951" athleteid="25199">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.97" eventid="5728" heatid="25717" lane="4" />
                <ENTRY entrytime="00:00:54.84" eventid="5744" heatid="25765" lane="5" />
                <ENTRY entrytime="00:02:10.00" eventid="1171" heatid="25820" lane="2" />
                <ENTRY entrytime="00:02:00.00" eventid="1195" heatid="25837" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lennart" gender="M" lastname="Köhler" nation="GER" license="354874" athleteid="25204">
              <ENTRIES>
                <ENTRY entrytime="00:02:23.85" eventid="1177" heatid="25664" lane="4" />
                <ENTRY entrytime="00:01:26.54" eventid="1141" heatid="25734" lane="2" />
                <ENTRY entrytime="00:00:31.76" eventid="5740" heatid="25760" lane="5" />
                <ENTRY entrytime="00:01:16.16" eventid="7773" heatid="25784" lane="4" />
                <ENTRY entrytime="00:01:14.64" eventid="1165" heatid="25819" lane="3" />
                <ENTRY entrytime="00:01:07.82" eventid="1189" heatid="25835" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Madlen" gender="F" lastname="Köthe" nation="GER" license="393115" athleteid="25211">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.40" eventid="5712" heatid="25688" lane="1" />
                <ENTRY entrytime="00:00:47.12" eventid="5744" heatid="25768" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="7788" heatid="25789" lane="2" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25802" lane="5" />
                <ENTRY entrytime="00:01:39.55" eventid="1195" heatid="25840" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Nadine" gender="F" lastname="Köttschau" nation="GER" license="392886" athleteid="25217">
              <ENTRIES>
                <ENTRY entrytime="00:03:41.42" eventid="1183" heatid="25667" lane="6" />
                <ENTRY entrytime="00:00:46.11" eventid="5728" heatid="25725" lane="6" />
                <ENTRY entrytime="00:02:00.63" eventid="1135" heatid="25738" lane="1" />
                <ENTRY entrytime="00:01:48.73" eventid="7788" heatid="25789" lane="4" />
                <ENTRY entrytime="00:01:44.97" eventid="1171" heatid="25822" lane="5" />
                <ENTRY entrytime="00:01:33.88" eventid="1195" heatid="25842" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Nina" gender="F" lastname="Köttschau" nation="GER" license="392885" athleteid="25224">
              <ENTRIES>
                <ENTRY entrytime="00:03:35.22" eventid="1183" heatid="25667" lane="4" />
                <ENTRY entrytime="00:00:46.05" eventid="5728" heatid="25725" lane="1" />
                <ENTRY entrytime="00:01:51.72" eventid="1135" heatid="25741" lane="2" />
                <ENTRY entrytime="00:00:42.13" eventid="1123" heatid="25815" lane="1" />
                <ENTRY entrytime="00:01:43.96" eventid="1171" heatid="25822" lane="2" />
                <ENTRY entrytime="00:01:32.61" eventid="1195" heatid="25842" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Paolo Emanuele" gender="M" lastname="Marzo" nation="GER" license="420810" athleteid="25237">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.30" eventid="5702" heatid="25676" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5724" heatid="25707" lane="6" />
                <ENTRY entrytime="00:01:07.69" eventid="5740" heatid="25747" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Julina" gender="F" lastname="Michel" nation="GER" license="404917" athleteid="25241">
              <ENTRIES>
                <ENTRY entrytime="00:03:16.03" eventid="1183" heatid="25670" lane="2" />
                <ENTRY entrytime="00:00:43.41" eventid="5728" heatid="25726" lane="3" />
                <ENTRY entrytime="00:00:37.35" eventid="5744" heatid="25775" lane="2" />
                <ENTRY entrytime="00:01:48.11" eventid="7788" heatid="25789" lane="3" />
                <ENTRY entrytime="00:01:29.59" eventid="1171" heatid="25824" lane="5" />
                <ENTRY entrytime="00:01:29.56" eventid="1195" heatid="25844" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Emilia" gender="F" lastname="Miller" nation="GER" license="414883" athleteid="25248">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.50" eventid="5712" heatid="25689" lane="1" />
                <ENTRY entrytime="00:00:55.78" eventid="5728" heatid="25720" lane="4" />
                <ENTRY entrytime="00:00:51.06" eventid="5744" heatid="25766" lane="6" />
                <ENTRY entrytime="00:00:30.00" eventid="7809" heatid="25799" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Fabian" gender="M" lastname="Muschik" nation="GER" license="373922" athleteid="25253">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.65" eventid="1177" heatid="25664" lane="3" />
                <ENTRY entrytime="00:00:37.10" eventid="5702" heatid="25684" lane="3" />
                <ENTRY entrytime="00:01:20.56" eventid="1141" heatid="25734" lane="3" />
                <ENTRY entrytime="00:00:29.72" eventid="5740" heatid="25760" lane="4" />
                <ENTRY entrytime="00:01:14.53" eventid="7773" heatid="25784" lane="3" />
                <ENTRY entrytime="00:01:06.15" eventid="1189" heatid="25835" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lia" gender="F" lastname="Puzicha" nation="GER" license="390447" athleteid="25260">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.88" eventid="5712" heatid="25696" lane="1" />
                <ENTRY entrytime="00:00:51.22" eventid="5728" heatid="25722" lane="2" />
                <ENTRY entrytime="00:01:55.07" eventid="1135" heatid="25740" lane="5" />
                <ENTRY entrytime="00:01:44.92" eventid="7788" heatid="25790" lane="2" />
                <ENTRY entrytime="00:01:50.54" eventid="1171" heatid="25821" lane="4" />
                <ENTRY entrytime="00:01:40.02" eventid="1195" heatid="25840" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Adrian" gender="M" lastname="Rohn" nation="GER" license="390446" athleteid="25267">
              <ENTRIES>
                <ENTRY entrytime="00:02:59.76" eventid="1177" heatid="25663" lane="1" />
                <ENTRY entrytime="00:00:44.67" eventid="5724" heatid="25714" lane="6" />
                <ENTRY entrytime="00:01:35.69" eventid="7773" heatid="25783" lane="6" />
                <ENTRY entrytime="00:01:34.06" eventid="1165" heatid="25818" lane="2" />
                <ENTRY entrytime="00:01:23.86" eventid="1189" heatid="25833" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Pierre" gender="M" lastname="Rudat" nation="GER" license="406826" athleteid="25273">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.44" eventid="5702" heatid="25674" lane="4" />
                <ENTRY entrytime="00:01:04.34" eventid="5724" heatid="25706" lane="1" />
                <ENTRY entrytime="00:00:49.25" eventid="5740" heatid="25751" lane="4" />
                <ENTRY entrytime="00:02:15.00" eventid="7773" heatid="25779" lane="1" />
                <ENTRY entrytime="00:01:10.00" eventid="1117" heatid="25804" lane="2" />
                <ENTRY entrytime="00:01:57.65" eventid="1189" heatid="25827" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Artur" gender="M" lastname="Schmal" nation="GER" license="425765" athleteid="25280">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.03" eventid="5702" heatid="25674" lane="1" />
                <ENTRY entrytime="00:01:06.50" eventid="5724" heatid="25705" lane="5" />
                <ENTRY entrytime="00:00:57.12" eventid="5740" heatid="25750" lane="6" />
                <ENTRY entrytime="00:00:35.00" eventid="7804" heatid="25795" lane="1" />
                <ENTRY entrytime="00:02:07.00" eventid="1189" heatid="25826" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Sophie" gender="F" lastname="Schmidt" nation="GER" license="420809" athleteid="25286">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25687" lane="5" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25716" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25763" lane="1" />
                <ENTRY entrytime="00:02:10.00" eventid="1195" heatid="25836" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leanora" gender="F" lastname="Sebeld" nation="GER" license="414884" athleteid="25291">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.44" eventid="5712" heatid="25689" lane="2" />
                <ENTRY entrytime="00:00:46.88" eventid="5728" heatid="25724" lane="5" />
                <ENTRY entrytime="00:00:38.10" eventid="5744" heatid="25774" lane="2" />
                <ENTRY entrytime="00:01:46.65" eventid="1171" heatid="25821" lane="3" />
                <ENTRY entrytime="00:01:30.16" eventid="1195" heatid="25843" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Veit-Josef" gender="M" lastname="Seidel" nation="GER" license="393117" athleteid="25297">
              <ENTRIES>
                <ENTRY entrytime="00:03:26.43" eventid="1177" heatid="25661" lane="6" />
                <ENTRY entrytime="00:00:47.15" eventid="5724" heatid="25712" lane="3" />
                <ENTRY entrytime="00:00:38.21" eventid="5740" heatid="25757" lane="5" />
                <ENTRY entrytime="00:01:37.06" eventid="7773" heatid="25782" lane="4" />
                <ENTRY entrytime="00:01:28.57" eventid="1189" heatid="25831" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Marc Steven" gender="M" lastname="Smirnov" nation="GER" license="417321" athleteid="25303">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.03" eventid="5702" heatid="25675" lane="2" />
                <ENTRY entrytime="00:00:57.06" eventid="5724" heatid="25708" lane="2" />
                <ENTRY entrytime="00:00:49.32" eventid="5740" heatid="25751" lane="2" />
                <ENTRY entrytime="00:02:15.00" eventid="7773" heatid="25779" lane="6" />
                <ENTRY entrytime="00:01:10.00" eventid="1117" heatid="25804" lane="4" />
                <ENTRY entrytime="00:01:57.94" eventid="1189" heatid="25826" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Elisabeth" gender="F" lastname="Strecker" nation="GER" license="406754" athleteid="25310">
              <ENTRIES>
                <ENTRY entrytime="00:03:19.87" eventid="1183" heatid="25670" lane="6" />
                <ENTRY entrytime="00:00:44.78" eventid="5728" heatid="25726" lane="5" />
                <ENTRY entrytime="00:00:39.41" eventid="5744" heatid="25773" lane="5" />
                <ENTRY entrytime="00:00:47.53" eventid="1123" heatid="25813" lane="2" />
                <ENTRY entrytime="00:01:36.81" eventid="1171" heatid="25823" lane="2" />
                <ENTRY entrytime="00:01:29.42" eventid="1195" heatid="25844" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Mark" gender="M" lastname="Sukhov" nation="GER" license="406821" athleteid="25317">
              <ENTRIES>
                <ENTRY entrytime="00:03:01.65" eventid="1177" heatid="25662" lane="3" />
                <ENTRY entrytime="00:01:45.00" eventid="1103" heatid="25699" lane="2" />
                <ENTRY entrytime="00:00:37.40" eventid="5740" heatid="25757" lane="3" />
                <ENTRY entrytime="00:01:34.02" eventid="1165" heatid="25818" lane="4" />
                <ENTRY entrytime="00:03:20.00" eventid="5655" heatid="25849" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Robin" gender="M" lastname="Tiede" nation="GER" license="404730" athleteid="25323">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.62" eventid="5702" heatid="25681" lane="6" />
                <ENTRY entrytime="00:00:45.48" eventid="5724" heatid="25713" lane="4" />
                <ENTRY entrytime="00:00:41.65" eventid="5740" heatid="25755" lane="5" />
                <ENTRY entrytime="00:01:40.00" eventid="7773" heatid="25782" lane="6" />
                <ENTRY entrytime="00:01:41.47" eventid="1165" heatid="25817" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Corali" gender="F" lastname="Walther" nation="GER" license="0" athleteid="25329">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.00" eventid="5664" heatid="25617" lane="4" />
                <ENTRY entrytime="00:00:25.00" eventid="5682" heatid="25631" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="7696" heatid="25638" lane="1" />
                <ENTRY entrytime="00:00:40.00" eventid="5690" heatid="25645" lane="4" />
                <ENTRY entrytime="00:00:35.00" eventid="5698" heatid="25655" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Mara Malin" gender="F" lastname="Walther" nation="GER" license="362627" athleteid="25335">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.36" eventid="5712" heatid="25697" lane="1" />
                <ENTRY entrytime="00:01:48.80" eventid="1135" heatid="25743" lane="6" />
                <ENTRY entrytime="00:00:39.58" eventid="5744" heatid="25773" lane="1" />
                <ENTRY entrytime="00:00:50.67" eventid="1123" heatid="25811" lane="2" />
                <ENTRY entrytime="00:01:40.17" eventid="1171" heatid="25823" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Helena" gender="F" lastname="Willared" nation="GER" license="368438" athleteid="25341">
              <ENTRIES>
                <ENTRY entrytime="00:03:24.14" eventid="1183" heatid="25669" lane="1" />
                <ENTRY entrytime="00:01:49.36" eventid="1135" heatid="25742" lane="2" />
                <ENTRY entrytime="00:00:37.97" eventid="5744" heatid="25774" lane="3" />
                <ENTRY entrytime="00:01:41.39" eventid="7788" heatid="25791" lane="6" />
                <ENTRY entrytime="00:01:40.70" eventid="1171" heatid="25822" lane="3" />
                <ENTRY entrytime="00:01:29.42" eventid="1195" heatid="25844" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6621" nation="GER" region="02" clubid="24230" name="SG Rödental">
          <ATHLETES>
            <ATHLETE birthdate="2010-01-01" firstname="Esther" gender="F" lastname="Amberg" nation="GER" license="420966" athleteid="24231">
              <ENTRIES>
                <ENTRY entrytime="00:03:55.00" eventid="1183" heatid="25666" lane="1" />
                <ENTRY entrytime="00:00:55.62" eventid="5728" heatid="25721" lane="6" />
                <ENTRY entrytime="00:02:04.51" eventid="7788" heatid="25786" lane="4" />
                <ENTRY entrytime="00:00:32.00" eventid="7809" heatid="25799" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Theresa" gender="F" lastname="Dressel" nation="GER" license="0" athleteid="24236">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.00" eventid="5664" heatid="25616" lane="5" />
                <ENTRY entrytime="00:00:43.00" eventid="5682" heatid="25629" lane="1" />
                <ENTRY entrytime="00:00:39.00" eventid="5690" heatid="25645" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="25653" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Hannes" gender="M" lastname="Endruweit" nation="GER" license="0" athleteid="24241">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="1053" heatid="25610" lane="6" />
                <ENTRY entrytime="00:00:35.00" eventid="5678" heatid="25624" lane="1" />
                <ENTRY entrytime="00:00:35.00" eventid="7691" heatid="25634" lane="4" />
                <ENTRY entrytime="00:00:55.00" eventid="7701" heatid="25657" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Jannik" gender="M" lastname="Endruweit" nation="GER" license="380996" athleteid="24246">
              <ENTRIES>
                <ENTRY entrytime="00:02:48.61" eventid="1177" heatid="25663" lane="3" />
                <ENTRY entrytime="00:01:29.55" eventid="1103" heatid="25700" lane="5" />
                <ENTRY entrytime="00:01:27.58" eventid="7773" heatid="25783" lane="3" />
                <ENTRY entrytime="00:00:18.00" eventid="7804" heatid="25797" lane="3" />
                <ENTRY entrytime="00:01:15.20" eventid="1189" heatid="25834" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Emely" gender="F" lastname="Gräser" nation="GER" license="367553" athleteid="24252">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.42" eventid="5728" heatid="25727" lane="3" />
                <ENTRY entrytime="00:00:34.05" eventid="5744" heatid="25776" lane="3" />
                <ENTRY entrytime="00:01:28.86" eventid="7788" heatid="25793" lane="4" />
                <ENTRY entrytime="00:01:23.08" eventid="1171" heatid="25824" lane="3" />
                <ENTRY entrytime="00:01:14.45" eventid="1195" heatid="25847" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Till" gender="M" lastname="Gräser" nation="GER" license="404231" athleteid="24258">
              <ENTRIES>
                <ENTRY entrytime="00:03:36.42" eventid="1177" heatid="25660" lane="2" />
                <ENTRY entrytime="00:00:48.88" eventid="5724" heatid="25711" lane="3" />
                <ENTRY entrytime="00:00:38.51" eventid="5740" heatid="25757" lane="1" />
                <ENTRY entrytime="00:00:30.00" eventid="7804" heatid="25795" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Anne-Lotte" gender="F" lastname="Hofbauer" nation="GER" license="417943" athleteid="24263">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.70" eventid="5712" heatid="25690" lane="6" />
                <ENTRY entrytime="00:02:19.64" eventid="1135" heatid="25735" lane="3" />
                <ENTRY entrytime="00:00:47.02" eventid="5744" heatid="25769" lane="6" />
                <ENTRY entrytime="00:02:10.00" eventid="1171" heatid="25820" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lennart" gender="M" lastname="Hofbauer" nation="GER" license="364856" athleteid="24268">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.44" eventid="5702" heatid="25684" lane="1" />
                <ENTRY entrytime="00:00:46.66" eventid="5724" heatid="25713" lane="1" />
                <ENTRY entrytime="00:00:33.97" eventid="5740" heatid="25759" lane="4" />
                <ENTRY entrytime="00:01:33.00" eventid="7773" heatid="25783" lane="5" />
                <ENTRY entrytime="00:01:14.96" eventid="1189" heatid="25834" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Jonathan" gender="M" lastname="Kohles" nation="GER" license="373339" athleteid="24274">
              <ENTRIES>
                <ENTRY entrytime="00:01:30.83" eventid="1103" heatid="25700" lane="1" />
                <ENTRY entrytime="00:01:23.99" eventid="1141" heatid="25734" lane="4" />
                <ENTRY entrytime="00:01:22.00" eventid="7773" heatid="25784" lane="5" />
                <ENTRY entrytime="00:00:37.00" eventid="1117" heatid="25808" lane="4" />
                <ENTRY entrytime="00:01:13.89" eventid="1189" heatid="25834" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Sophia" gender="F" lastname="Lamik" nation="GER" license="0" athleteid="24280">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.00" eventid="5664" heatid="25614" lane="2" />
                <ENTRY entrytime="00:00:42.00" eventid="7696" heatid="25638" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="25653" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="7706" heatid="25658" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Arne" gender="M" lastname="Mesch" nation="GER" license="361790" athleteid="24285">
              <ENTRIES>
                <ENTRY entrytime="00:02:33.29" eventid="1177" heatid="25664" lane="1" />
                <ENTRY entrytime="00:00:37.81" eventid="5724" heatid="25714" lane="4" />
                <ENTRY entrytime="00:01:19.61" eventid="7773" heatid="25784" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="1117" heatid="25808" lane="2" />
                <ENTRY entrytime="00:01:08.15" eventid="1189" heatid="25835" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Tobais Damian" gender="M" lastname="Schiebert" nation="GER" license="429408" athleteid="24291">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5702" heatid="25674" lane="2" />
                <ENTRY entrytime="00:01:10.00" eventid="5724" heatid="25704" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="25748" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Manuel" gender="M" lastname="Staffel" nation="GER" license="364847" athleteid="24295">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.41" eventid="1177" heatid="25663" lane="2" />
                <ENTRY entrytime="00:00:35.54" eventid="5740" heatid="25758" lane="3" />
                <ENTRY entrytime="00:01:38.64" eventid="7773" heatid="25782" lane="1" />
                <ENTRY entrytime="00:01:38.02" eventid="1165" heatid="25818" lane="5" />
                <ENTRY entrytime="00:01:17.76" eventid="1189" heatid="25834" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Istvan" gender="M" lastname="Sziklavari" nation="GER" license="000000" athleteid="25433">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5702" heatid="25673" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2014-01-01" firstname="Nandor" gender="M" lastname="Sziklavari" nation="GER" license="000000" athleteid="25431">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25607" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lea" gender="F" lastname="Tarrach" nation="GER" license="373337" athleteid="24301">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.25" eventid="5712" heatid="25698" lane="4" />
                <ENTRY entrytime="00:01:34.79" eventid="1135" heatid="25745" lane="4" />
                <ENTRY entrytime="00:00:36.21" eventid="5744" heatid="25776" lane="6" />
                <ENTRY entrytime="00:01:38.00" eventid="7788" heatid="25791" lane="5" />
                <ENTRY entrytime="00:01:21.11" eventid="1195" heatid="25846" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lina" gender="F" lastname="Tarrach" nation="GER" license="417942" athleteid="24307">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.39" eventid="5712" heatid="25692" lane="4" />
                <ENTRY entrytime="00:01:02.40" eventid="5728" heatid="25717" lane="5" />
                <ENTRY entrytime="00:02:07.72" eventid="1135" heatid="25737" lane="6" />
                <ENTRY entrytime="00:02:05.00" eventid="1195" heatid="25837" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Johanna" gender="F" lastname="Thiem" nation="GER" license="404230" athleteid="24312">
              <ENTRIES>
                <ENTRY entrytime="00:03:33.93" eventid="1183" heatid="25668" lane="6" />
                <ENTRY entrytime="00:01:59.86" eventid="7788" heatid="25787" lane="3" />
                <ENTRY entrytime="00:00:50.56" eventid="1123" heatid="25811" lane="4" />
                <ENTRY entrytime="00:01:48.13" eventid="1195" heatid="25839" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Vanessa" gender="F" lastname="Thiem" nation="GER" license="404232" athleteid="24317">
              <ENTRIES>
                <ENTRY entrytime="00:02:57.28" eventid="1183" heatid="25672" lane="1" />
                <ENTRY entrytime="00:00:35.95" eventid="5744" heatid="25776" lane="2" />
                <ENTRY entrytime="00:01:34.05" eventid="7788" heatid="25792" lane="5" />
                <ENTRY entrytime="00:00:42.81" eventid="1123" heatid="25815" lane="6" />
                <ENTRY entrytime="00:01:19.53" eventid="1195" heatid="25847" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Alina" gender="F" lastname="Zeder" nation="GER" license="0" athleteid="24323">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.00" eventid="5664" heatid="25614" lane="3" />
                <ENTRY entrytime="00:00:39.00" eventid="7696" heatid="25638" lane="5" />
                <ENTRY entrytime="00:00:37.00" eventid="5690" heatid="25646" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="25653" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Bastian" gender="M" lastname="Zetzmann" nation="GER" license="392527" athleteid="24328">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.55" eventid="5702" heatid="25680" lane="5" />
                <ENTRY entrytime="00:02:00.73" eventid="1141" heatid="25730" lane="4" />
                <ENTRY entrytime="00:02:05.00" eventid="7773" heatid="25779" lane="2" />
                <ENTRY entrytime="00:01:48.00" eventid="1189" heatid="25828" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6655" nation="GER" region="02" clubid="24810" name="TSG Nürnberg">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="Leni" gender="F" lastname="Amadasun" nation="GER" license="407651" athleteid="25488">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.25" eventid="5712" heatid="25694" lane="5" />
                <ENTRY entrytime="00:01:55.00" eventid="1135" heatid="25740" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="7788" heatid="25789" lane="1" />
                <ENTRY entrytime="00:00:47.63" eventid="1123" heatid="25813" lane="1" />
                <ENTRY entrytime="00:01:38.09" eventid="1195" heatid="25841" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Alexey" gender="M" lastname="Antonkin" nation="GER" license="392619" athleteid="25494">
              <ENTRIES>
                <ENTRY entrytime="00:03:12.58" eventid="1177" heatid="25662" lane="6" />
                <ENTRY entrytime="00:00:46.45" eventid="5724" heatid="25713" lane="2" />
                <ENTRY entrytime="00:00:36.52" eventid="5740" heatid="25758" lane="2" />
                <ENTRY entrytime="00:00:55.47" eventid="1117" heatid="25805" lane="5" />
                <ENTRY entrytime="00:01:45.00" eventid="1165" heatid="25817" lane="5" />
                <ENTRY entrytime="00:01:26.00" eventid="1189" heatid="25832" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Alexander" gender="M" lastname="Eisler" nation="GER" license="0" athleteid="25573">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1177" heatid="25659" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5724" heatid="25707" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="5740" heatid="25750" lane="4" />
                <ENTRY entrytime="NT" eventid="1117" heatid="25804" lane="5" />
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25828" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Stas" gender="M" lastname="Eisler" nation="GER" license="0" athleteid="25579">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.00" eventid="5702" heatid="25682" lane="4" />
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25730" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="5740" heatid="25751" lane="1" />
                <ENTRY entrytime="00:00:25.00" eventid="7804" heatid="25797" lane="1" />
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25828" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Laura" gender="F" lastname="Evseenkov" nation="GER" license="404373" athleteid="25501">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.45" eventid="5712" heatid="25693" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="25738" lane="3" />
                <ENTRY entrytime="00:01:57.24" eventid="7788" heatid="25788" lane="6" />
                <ENTRY entrytime="00:00:30.00" eventid="7809" heatid="25800" lane="5" />
                <ENTRY entrytime="00:01:51.13" eventid="1195" heatid="25839" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Kim" gender="F" lastname="Forster" nation="GER" license="330020" athleteid="24811">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.02" eventid="5712" heatid="25698" lane="3" />
                <ENTRY entrytime="00:01:37.67" eventid="1135" heatid="25745" lane="5" />
                <ENTRY entrytime="00:01:33.64" eventid="7788" heatid="25792" lane="2" />
                <ENTRY entrytime="00:01:34.17" eventid="1171" heatid="25823" lane="4" />
                <ENTRY entrytime="00:01:23.70" eventid="1195" heatid="25845" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Sandrine" gender="F" lastname="Fuchs" nation="GER" license="407650" athleteid="25507">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25718" lane="3" />
                <ENTRY entrytime="00:00:59.97" eventid="5744" heatid="25763" lane="2" />
                <ENTRY entrytime="00:02:00.00" eventid="7788" heatid="25787" lane="4" />
                <ENTRY entrytime="00:00:30.00" eventid="7809" heatid="25800" lane="2" />
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25687" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Michael" gender="M" lastname="Geng" nation="GER" license="0" athleteid="25567">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="5702" heatid="25679" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25731" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5740" heatid="25750" lane="2" />
                <ENTRY entrytime="00:00:30.00" eventid="7804" heatid="25795" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="1165" heatid="25817" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lorena" gender="F" lastname="Graz" nation="GER" license="392620" athleteid="25513">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.51" eventid="5712" heatid="25697" lane="6" />
                <ENTRY entrytime="00:01:51.80" eventid="1135" heatid="25741" lane="5" />
                <ENTRY entrytime="00:00:42.06" eventid="5744" heatid="25771" lane="6" />
                <ENTRY entrytime="00:01:55.00" eventid="1171" heatid="25821" lane="1" />
                <ENTRY entrytime="00:01:41.06" eventid="1195" heatid="25840" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lorin" gender="F" lastname="Karakas" nation="GER" license="000000" athleteid="25600">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5712" heatid="25690" lane="2" />
                <ENTRY entrytime="00:00:30.00" eventid="7809" heatid="25800" lane="6" />
                <ENTRY entrytime="00:02:00.00" eventid="7788" heatid="25787" lane="5" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="25764" lane="4" />
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="25738" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lawan" gender="M" lastname="Karwan Farik" nation="GER" license="393140" athleteid="25868">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="5702" heatid="25679" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5724" heatid="25706" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25731" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="25748" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="7804" heatid="25795" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Anna" gender="F" lastname="Kießling" nation="GER" license="417716" athleteid="25519">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5712" heatid="25690" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="25738" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="5744" heatid="25766" lane="5" />
                <ENTRY entrytime="00:01:50.00" eventid="7788" heatid="25789" lane="5" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25802" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Valeria Alexandra" gender="F" lastname="Nekrasov" nation="GER" license="392621" athleteid="25525">
              <ENTRIES>
                <ENTRY entrytime="00:01:40.00" eventid="1111" heatid="25703" lane="1" />
                <ENTRY entrytime="00:01:36.77" eventid="1135" heatid="25745" lane="2" />
                <ENTRY entrytime="00:01:35.09" eventid="7788" heatid="25791" lane="3" />
                <ENTRY entrytime="00:00:41.48" eventid="1123" heatid="25815" lane="2" />
                <ENTRY entrytime="00:01:25.33" eventid="1171" heatid="25824" lane="2" />
                <ENTRY entrytime="00:04:00.00" eventid="5661" heatid="25850" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Jurij" gender="M" lastname="Pandeleer" nation="GER" license="0" athleteid="25595">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5702" heatid="25677" lane="5" />
                <ENTRY entrytime="NT" eventid="5724" heatid="25704" lane="6" />
                <ENTRY entrytime="NT" eventid="1141" heatid="25729" lane="6" />
                <ENTRY entrytime="NT" eventid="5740" heatid="25746" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Elisa" gender="F" lastname="Peter" nation="GER" license="0" athleteid="25585">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5712" heatid="25690" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25719" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="5744" heatid="25766" lane="4" />
                <ENTRY entrytime="00:00:30.00" eventid="7809" heatid="25799" lane="4" />
                <ENTRY entrytime="00:01:55.00" eventid="1195" heatid="25838" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Tobias" gender="M" lastname="Rhau" nation="GER" license="421150" athleteid="25532">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.55" eventid="5702" heatid="25678" lane="2" />
                <ENTRY entrytime="00:00:49.91" eventid="5740" heatid="25751" lane="5" />
                <ENTRY entrytime="00:01:55.00" eventid="7773" heatid="25780" lane="5" />
                <ENTRY entrytime="NT" eventid="1117" heatid="25804" lane="1" />
                <ENTRY entrytime="00:01:57.38" eventid="1189" heatid="25827" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Leila" gender="F" lastname="Schomleu" nation="GER" license="0" athleteid="25538">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.00" eventid="5664" heatid="25615" lane="2" />
                <ENTRY entrytime="00:00:45.00" eventid="5682" heatid="25628" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="25644" lane="1" />
                <ENTRY entrytime="00:00:46.00" eventid="5698" heatid="25654" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Tamina" gender="F" lastname="Schomleu" nation="GER" license="0" athleteid="25543">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.00" eventid="5664" heatid="25615" lane="6" />
                <ENTRY entrytime="00:00:45.00" eventid="5682" heatid="25628" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25636" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5690" heatid="25644" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="5698" heatid="25653" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lena" gender="F" lastname="Schreiber" nation="GER" license="392618" athleteid="25549">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.18" eventid="5712" heatid="25694" lane="2" />
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="25739" lane="6" />
                <ENTRY entrytime="00:02:00.00" eventid="7788" heatid="25787" lane="2" />
                <ENTRY entrytime="00:00:30.00" eventid="1123" heatid="25815" lane="3" />
                <ENTRY entrytime="00:01:50.18" eventid="1195" heatid="25839" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Jakob" gender="M" lastname="Sickmüller" nation="GER" license="359484" athleteid="25555">
              <ENTRIES>
                <ENTRY entrytime="00:03:30.00" eventid="1177" heatid="25660" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="1141" heatid="25732" lane="1" />
                <ENTRY entrytime="00:01:50.00" eventid="7773" heatid="25780" lane="3" />
                <ENTRY entrytime="00:01:34.74" eventid="1189" heatid="25830" lane="2" />
                <ENTRY entrytime="00:03:50.00" eventid="5655" heatid="25848" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Gleb" gender="M" lastname="Welsch" nation="GER" license="000000" athleteid="25852">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5702" heatid="25677" lane="2" />
                <ENTRY entrytime="00:20:00.00" eventid="1141" heatid="25729" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="5740" heatid="25750" lane="3" />
                <ENTRY entrytime="00:00:30.00" eventid="7804" heatid="25796" lane="6" />
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25827" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4502" nation="GER" region="02" clubid="24023" name="TSV Zirndorf">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Jana" gender="F" lastname="Ammon" nation="GER" license="398728" athleteid="24024">
              <ENTRIES>
                <ENTRY entrytime="00:03:00.00" eventid="1183" heatid="25671" lane="3" />
                <ENTRY entrytime="00:01:40.00" eventid="1111" heatid="25703" lane="5" />
                <ENTRY entrytime="00:00:41.63" eventid="5744" heatid="25771" lane="1" />
                <ENTRY entrytime="00:01:46.09" eventid="1171" heatid="25822" lane="1" />
                <ENTRY entrytime="00:01:27.68" eventid="1195" heatid="25844" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Marco" gender="M" lastname="Ammon" nation="GER" license="398727" athleteid="24030">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.00" eventid="1177" heatid="25663" lane="4" />
                <ENTRY entrytime="00:01:48.15" eventid="1141" heatid="25732" lane="5" />
                <ENTRY entrytime="00:01:38.56" eventid="7773" heatid="25782" lane="5" />
                <ENTRY entrytime="00:00:46.85" eventid="1117" heatid="25807" lane="2" />
                <ENTRY entrytime="00:02:50.00" eventid="5655" heatid="25849" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Alissa" gender="F" lastname="Bader" nation="GER" license="428030" athleteid="24036">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.00" eventid="1183" heatid="25671" lane="1" />
                <ENTRY entrytime="00:00:50.28" eventid="5712" heatid="25697" lane="5" />
                <ENTRY entrytime="00:01:56.25" eventid="1135" heatid="25740" lane="6" />
                <ENTRY entrytime="00:00:40.06" eventid="5744" heatid="25772" lane="2" />
                <ENTRY entrytime="00:01:36.53" eventid="1195" heatid="25841" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Mia" gender="F" lastname="Großhauser" nation="GER" license="420483" athleteid="24042">
              <ENTRIES>
                <ENTRY entrytime="00:03:10.00" eventid="1183" heatid="25671" lane="6" />
                <ENTRY entrytime="00:01:59.09" eventid="1135" heatid="25739" lane="1" />
                <ENTRY entrytime="00:01:53.94" eventid="7788" heatid="25788" lane="5" />
                <ENTRY entrytime="00:00:25.12" eventid="7809" heatid="25801" lane="5" />
                <ENTRY entrytime="00:01:35.78" eventid="1195" heatid="25841" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Josefine" gender="F" lastname="Mendler" nation="GER" license="420484" athleteid="24048">
              <ENTRIES>
                <ENTRY entrytime="00:03:40.00" eventid="1183" heatid="25667" lane="1" />
                <ENTRY entrytime="00:01:08.35" eventid="5728" heatid="25716" lane="2" />
                <ENTRY entrytime="00:02:08.52" eventid="1135" heatid="25736" lane="3" />
                <ENTRY entrytime="00:02:05.00" eventid="7788" heatid="25786" lane="2" />
                <ENTRY entrytime="00:02:02.26" eventid="1195" heatid="25837" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Simona" gender="F" lastname="Paschold" nation="GER" license="398731" athleteid="24054">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.74" eventid="1183" heatid="25672" lane="4" />
                <ENTRY entrytime="00:00:45.09" eventid="5728" heatid="25725" lane="4" />
                <ENTRY entrytime="00:01:37.69" eventid="1135" heatid="25745" lane="1" />
                <ENTRY entrytime="00:01:30.12" eventid="7788" heatid="25793" lane="1" />
                <ENTRY entrytime="00:00:45.56" eventid="1123" heatid="25814" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Tim Simon" gender="M" lastname="Paschold" nation="GER" license="428031" athleteid="24060">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.50" eventid="5702" heatid="25676" lane="5" />
                <ENTRY entrytime="00:01:05.93" eventid="5724" heatid="25705" lane="2" />
                <ENTRY entrytime="00:02:14.09" eventid="1141" heatid="25729" lane="4" />
                <ENTRY entrytime="00:00:48.87" eventid="5740" heatid="25752" lane="6" />
                <ENTRY entrytime="00:02:00.56" eventid="1189" heatid="25826" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
