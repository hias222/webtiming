<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SG Fürth" version="11.61084">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Fürth" name="42. Fürther Kinderschwimmen" course="SCM" deadline="2018-11-04" hostclub="SG Fürth" hostclub.url="http://www.sgfuerth.de" organizer="SG Fürth" organizer.url="http://www.sgfuerth.de" reservecount="2" startmethod="1" timing="AUTOMATIC" state="BY" nation="GER">
      <AGEDATE value="2018-11-10" type="YEAR" />
      <POOL name="Hallebad am Scherbsgraben" lanemin="1" lanemax="6" />
      <FACILITY city="Fürth" name="Hallebad am Scherbsgraben" nation="GER" state="BY" street="Scherbsgraben 15" zip="90765" />
      <POINTTABLE pointtableid="3011" name="FINA Point Scoring" version="2018" />
      <CONTACT city="Fürth" email="meldungen@sgfuerth.de" name="Matthias Fuchs" phone="09118101172" street="Lavendelweg 47" zip="90768" />
      <SESSIONS>
        <SESSION date="2018-11-10" daytime="08:30" endtime="10:56" number="1" officialmeeting="08:00" teamleadermeeting="08:15" warmupfrom="08:00" warmupuntil="08:25">
          <EVENTS>
            <EVENT eventid="5668" daytime="08:44" gender="M" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="103" name="25m Rückenbeine ohne Brett" stroke="UNKNOWN" code="25 Rub" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7651" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7652" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7653" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7654" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25756" daytime="08:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25757" daytime="08:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25758" daytime="08:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25759" daytime="08:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25760" daytime="08:48" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7691" daytime="09:06" gender="M" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="501" name="25m Kraulbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7692" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7693" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7694" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7695" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25774" daytime="09:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25775" daytime="09:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25776" daytime="09:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25777" daytime="09:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25778" daytime="09:12" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25779" daytime="09:14" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5678" daytime="08:58" gender="M" number="5" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7659" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7660" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7661" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7662" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25765" daytime="08:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25766" daytime="08:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25767" daytime="09:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25768" daytime="09:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25769" daytime="09:02" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7696" daytime="09:14" gender="F" number="8" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="501" name="25m Kraulbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7697" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7698" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7699" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7700" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25780" daytime="09:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25781" daytime="09:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25782" daytime="09:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25783" daytime="09:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25784" daytime="09:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25785" daytime="09:22" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7706" daytime="10:10" gender="F" number="14" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="502" name="25m Delphinbeine o. Brett" stroke="UNKNOWN" code="25 Dob" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7707" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7708" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7709" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7710" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25808" daytime="10:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25809" daytime="10:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5674" daytime="08:50" gender="F" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="103" name="25m Rückenbeine ohne Brett" stroke="UNKNOWN" code="25 Rub" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7655" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7656" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7657" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7658" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25761" daytime="08:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25762" daytime="08:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25763" daytime="08:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25764" daytime="08:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5686" daytime="09:44" gender="M" number="9" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="101" name="25m Brustbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7667" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7668" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7669" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7670" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25786" daytime="09:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25787" daytime="09:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25788" daytime="09:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25789" daytime="09:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25790" daytime="09:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25791" daytime="09:50" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5664" daytime="08:36" gender="F" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7647" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7648" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7649" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7650" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25750" daytime="08:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25751" daytime="08:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25752" daytime="08:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25753" daytime="08:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25754" daytime="08:42" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25755" daytime="08:42" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5682" daytime="09:02" gender="F" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7663" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7664" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7665" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7666" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25770" daytime="09:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25771" daytime="09:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25772" daytime="09:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25773" daytime="09:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5694" daytime="09:58" gender="M" number="11" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7675" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7676" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7677" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7678" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25797" daytime="09:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25798" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25799" daytime="10:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25800" daytime="10:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25801" daytime="10:04" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5690" daytime="09:52" gender="F" number="10" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="101" name="25m Brustbeine mit Brett" stroke="UNKNOWN" code="25 Frb" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7671" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7672" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7673" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7674" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25792" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25793" daytime="09:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25794" daytime="09:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25795" daytime="09:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25796" daytime="09:58" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5698" daytime="10:04" gender="F" number="12" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7679" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7680" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7681" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7682" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25802" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25803" daytime="10:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25804" daytime="10:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25805" daytime="10:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25806" daytime="10:08" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1053" daytime="08:30" gender="M" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7646" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="1055" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="1054" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="2915" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25744" daytime="08:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25745" daytime="08:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25746" daytime="08:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25747" daytime="08:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25748" daytime="08:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25749" daytime="08:36" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7701" daytime="10:10" gender="M" number="13" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" swimstyleid="502" name="25m Delphinbeine o. Brett" stroke="UNKNOWN" code="25 Dob" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7702" agemax="4" agemin="4" />
                <AGEGROUP agegroupid="7703" agemax="5" agemin="5" />
                <AGEGROUP agegroupid="7704" agemax="6" agemin="6" />
                <AGEGROUP agegroupid="7705" agemax="7" agemin="7" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25807" daytime="10:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="17217" role="REF" />
            <JUDGE number="2" officialid="26024" role="REF" />
            <JUDGE number="1" officialid="26026" role="STA" />
            <JUDGE number="2" officialid="26028" role="STA" />
            <JUDGE number="1" officialid="26030" role="ANN" />
            <JUDGE number="2" officialid="26032" role="ANN" />
            <JUDGE number="1" officialid="26034" role="AW" />
            <JUDGE number="2" officialid="17223" role="AW" />
            <JUDGE number="1" officialid="26037" role="CRS" />
            <JUDGE number="2" officialid="26039" role="CRS" />
            <JUDGE number="1" officialid="26041" role="JOS" />
            <JUDGE number="2" officialid="26043" role="JOS" />
            <JUDGE number="1" officialid="26045" role="CFIN" />
            <JUDGE number="1" officialid="26047" role="FIN" />
            <JUDGE number="2" officialid="26049" role="FIN" />
            <JUDGE number="1" officialid="26051" role="CTIK" />
            <JUDGE number="1" officialid="26053" role="TIK" />
            <JUDGE number="2" officialid="26055" role="TIK" />
            <JUDGE number="3" officialid="17185" role="TIK" />
            <JUDGE number="4" officialid="26058" role="TIK" />
            <JUDGE number="5" officialid="26060" role="TIK" />
            <JUDGE number="6" officialid="17212" role="TIK" />
            <JUDGE number="1" officialid="23676" role="RTIK" />
            <JUDGE number="1" officialid="26064" role="CIOT" />
            <JUDGE number="1" officialid="26066" role="IOT" />
            <JUDGE number="2" officialid="26068" role="IOT" />
          </JUDGES>
        </SESSION>
        <SESSION date="2018-11-10" daytime="12:00" endtime="19:12" number="2" officialmeeting="11:30" teamleadermeeting="11:30" warmupfrom="11:00" warmupuntil="11:55">
          <EVENTS>
            <EVENT eventid="7773" daytime="15:28" gender="M" number="27" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7781" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7782" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7783" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7784" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7785" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7786" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7787" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25929" daytime="15:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25930" daytime="15:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25931" daytime="15:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25932" daytime="15:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25933" daytime="15:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25934" daytime="15:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25935" daytime="15:42" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5744" daytime="15:06" gender="F" number="26" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23817" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23818" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23819" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23820" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23821" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23822" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23823" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25912" daytime="15:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25913" daytime="15:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25914" daytime="15:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25915" daytime="15:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25916" daytime="15:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25917" daytime="15:14" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25918" daytime="15:16" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25919" daytime="15:18" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25920" daytime="15:18" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25921" daytime="15:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25922" daytime="15:20" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25923" daytime="15:22" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="25924" daytime="15:22" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="25925" daytime="15:24" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="25926" daytime="15:24" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="25927" daytime="15:26" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="25928" daytime="15:26" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7809" daytime="16:44" gender="F" number="31" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7818" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7819" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7820" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7821" agemax="11" agemin="11" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25951" daytime="16:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25952" daytime="16:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25953" daytime="16:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25954" daytime="16:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25955" daytime="16:48" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="13:20" gender="M" number="19" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7721" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1105" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1104" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1107" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1106" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1109" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25848" daytime="13:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7788" daytime="15:44" gender="F" number="28" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7789" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7790" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7791" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7792" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7793" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7794" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7795" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25936" daytime="15:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25937" daytime="15:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25938" daytime="15:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25939" daytime="15:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25940" daytime="15:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25941" daytime="15:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25942" daytime="16:00" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25943" daytime="16:02" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25944" daytime="16:04" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25945" daytime="16:06" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="17:14" gender="F" number="35" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7837" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7838" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7839" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7840" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7841" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7842" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7843" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25973" daytime="17:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25974" daytime="17:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25975" daytime="17:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25976" daytime="17:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25977" daytime="17:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25978" daytime="17:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25979" daytime="17:28" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25980" daytime="17:30" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5702" daytime="12:46" gender="M" number="17" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23782" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23783" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23784" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23785" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23786" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23787" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23788" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25821" daytime="12:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25822" daytime="12:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25823" daytime="12:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25824" daytime="12:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25825" daytime="12:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25826" daytime="12:54" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25827" daytime="12:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25828" daytime="12:56" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25829" daytime="12:56" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25830" daytime="12:58" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25831" daytime="12:58" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25832" daytime="13:00" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5655" daytime="18:26" gender="M" number="38" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7870" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7871" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7872" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7873" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7874" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7875" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="26006" daytime="18:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="26007" daytime="18:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1177" daytime="12:00" gender="M" number="15" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7746" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7747" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7748" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7749" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7750" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7751" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25810" daytime="12:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25811" daytime="12:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25812" daytime="12:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25813" daytime="12:12" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5724" daytime="13:28" gender="M" number="21" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23796" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23797" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23798" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23799" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23800" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23801" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23802" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25852" daytime="13:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25853" daytime="13:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25854" daytime="13:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25855" daytime="13:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25856" daytime="13:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25857" daytime="13:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25858" daytime="13:38" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25859" daytime="13:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25860" daytime="13:40" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25861" daytime="13:42" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25862" daytime="13:42" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25863" daytime="13:44" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="17:58" gender="F" number="37" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7863" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7864" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7865" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7866" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7867" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7868" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7869" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25993" daytime="17:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25994" daytime="18:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25995" daytime="18:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25996" daytime="18:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25997" daytime="18:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25998" daytime="18:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25999" daytime="18:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="26000" daytime="18:14" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="26001" daytime="18:16" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="26002" daytime="18:18" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="26003" daytime="18:20" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="26004" daytime="18:22" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="26005" daytime="18:24" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5740" daytime="14:50" gender="M" number="25" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23810" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23811" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23812" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23813" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23814" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23815" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23816" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25898" daytime="14:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25899" daytime="14:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25900" daytime="14:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25901" daytime="14:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25902" daytime="14:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25903" daytime="14:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25904" daytime="14:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25905" daytime="15:00" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25906" daytime="15:02" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25907" daytime="15:02" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25908" daytime="15:04" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25909" daytime="15:04" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="25910" daytime="15:06" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="25911" daytime="15:06" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5661" daytime="18:34" gender="F" number="39" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7876" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7877" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7878" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7879" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7880" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7881" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="26008" daytime="18:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="26009" daytime="18:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="26010" daytime="18:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="26011" daytime="18:46" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="23774" daytime="16:08" gender="X" number="29" order="18" round="TIM" maxentries="1" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23775" agemax="14" agemin="8" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25946" daytime="16:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7804" daytime="16:40" gender="M" number="30" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7814" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7815" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7816" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7817" agemax="11" agemin="11" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25947" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25948" daytime="16:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25949" daytime="16:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25950" daytime="16:42" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5712" daytime="13:02" gender="F" number="18" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23789" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23790" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23791" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23792" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23793" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23794" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23795" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25833" daytime="13:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25834" daytime="13:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25835" daytime="13:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25836" daytime="13:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25837" daytime="13:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25838" daytime="13:08" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25839" daytime="13:10" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25840" daytime="13:12" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25841" daytime="13:12" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25842" daytime="13:14" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25843" daytime="13:14" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25844" daytime="13:16" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="25845" daytime="13:16" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="25846" daytime="13:18" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="25847" daytime="13:20" number="15" order="15" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" daytime="14:02" gender="M" number="23" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7759" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7760" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7761" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7762" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7763" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7764" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7765" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25878" daytime="14:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25879" daytime="14:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25880" daytime="14:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25881" daytime="14:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25882" daytime="14:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25883" daytime="14:16" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25884" daytime="14:18" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25885" daytime="14:20" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5728" daytime="13:44" gender="F" number="22" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23803" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23804" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23805" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23806" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23807" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23808" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23809" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25864" daytime="13:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25865" daytime="13:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25866" daytime="13:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25867" daytime="13:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25868" daytime="13:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25869" daytime="13:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25870" daytime="13:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25871" daytime="13:54" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25872" daytime="13:56" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25873" daytime="13:58" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25874" daytime="13:58" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25875" daytime="14:00" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="25876" daytime="14:00" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="25877" daytime="14:02" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="12:16" gender="F" number="16" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7753" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7754" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7755" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7756" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7757" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7758" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25814" daytime="12:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25815" daytime="12:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25816" daytime="12:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25817" daytime="12:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25818" daytime="12:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25819" daytime="12:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25820" daytime="12:42" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1189" daytime="17:32" gender="M" number="36" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7856" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7857" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7858" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7859" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7860" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7861" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7862" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25981" daytime="17:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25982" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25983" daytime="17:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25984" daytime="17:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25985" daytime="17:42" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25986" daytime="17:44" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25987" daytime="17:46" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25988" daytime="17:48" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25989" daytime="17:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25990" daytime="17:52" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25991" daytime="17:54" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25992" daytime="17:56" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="13:22" gender="F" number="20" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7722" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1112" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="1113" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1114" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="1115" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1116" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25849" daytime="13:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25850" daytime="13:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25851" daytime="13:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="14:22" gender="F" number="24" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7766" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7767" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7768" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7769" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7770" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7771" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7772" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25886" daytime="14:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25887" daytime="14:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25888" daytime="14:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25889" daytime="14:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25890" daytime="14:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25891" daytime="14:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="25892" daytime="14:38" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="25893" daytime="14:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="25894" daytime="14:42" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="25895" daytime="14:44" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="25896" daytime="14:46" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="25897" daytime="14:48" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="17:02" gender="M" number="34" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7830" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="7831" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="7832" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="7833" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="7834" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="7835" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="7836" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25967" daytime="17:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25968" daytime="17:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25969" daytime="17:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25970" daytime="17:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25971" daytime="17:12" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25972" daytime="17:14" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" daytime="16:48" gender="M" number="32" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23824" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23825" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23826" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23827" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23828" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23829" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23830" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25956" daytime="16:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25957" daytime="16:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25958" daytime="16:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25959" daytime="16:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25960" daytime="16:52" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1123" daytime="16:54" gender="F" number="33" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="450" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23831" agemax="8" agemin="8" />
                <AGEGROUP agegroupid="23832" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="23833" agemax="10" agemin="10" />
                <AGEGROUP agegroupid="23834" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="23835" agemax="12" agemin="12" />
                <AGEGROUP agegroupid="23836" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="23837" agemax="14" agemin="14" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="25961" daytime="16:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="25962" daytime="16:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="25963" daytime="16:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="25964" daytime="16:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="25965" daytime="17:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="25966" daytime="17:00" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE number="1" officialid="17217" role="REF" />
            <JUDGE number="2" officialid="17223" role="REF" />
            <JUDGE number="1" officialid="26026" role="STA" />
            <JUDGE number="2" officialid="26028" role="STA" />
            <JUDGE number="1" officialid="26030" role="ANN" />
            <JUDGE number="2" officialid="26032" role="ANN" />
            <JUDGE number="1" officialid="26034" role="AW" />
            <JUDGE number="1" officialid="26037" role="CRS" />
            <JUDGE number="2" officialid="26039" role="CRS" />
            <JUDGE number="1" officialid="26095" role="JOS" />
            <JUDGE number="2" officialid="26096" role="JOS" />
            <JUDGE number="1" officialid="26097" role="CFIN" />
            <JUDGE number="1" officialid="26098" role="FIN" />
            <JUDGE number="2" officialid="26099" role="FIN" />
            <JUDGE number="1" officialid="26100" role="CTIK" />
            <JUDGE number="1" officialid="26101" role="TIK" />
            <JUDGE number="2" officialid="26102" role="TIK" />
            <JUDGE number="3" officialid="17185" role="TIK" />
            <JUDGE number="4" officialid="17182" role="TIK" />
            <JUDGE number="5" officialid="26103" role="TIK" />
            <JUDGE number="6" officialid="17212" role="TIK" />
            <JUDGE number="1" officialid="26104" role="RTIK" />
            <JUDGE number="2" officialid="26060" role="RTIK" />
            <JUDGE number="11" officialid="26110" role="TIK" />
            <JUDGE number="12" officialid="23615" role="TIK" />
            <JUDGE number="13" officialid="26115" role="TIK" />
            <JUDGE number="14" officialid="26116" role="TIK" />
            <JUDGE number="15" officialid="26117" role="TIK" />
            <JUDGE number="16" officialid="26118" role="TIK" />
            <JUDGE number="1" officialid="23767" role="CIOT" />
            <JUDGE number="1" officialid="26106" role="IOT" />
            <JUDGE number="2" officialid="26107" role="IOT" />
          </JUDGES>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="4363" nation="GER" region="02" clubid="7967" name="1. SV Nördlingen" />
        <CLUB type="CLUB" code="4163" nation="GER" region="02" clubid="7942" name="1.FCN Schwimmen">
          <OFFICIALS>
            <OFFICIAL officialid="17214" firstname="Petra" gender="F" lastname="Forster" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4167" nation="GER" region="02" clubid="7902" name="1.SC Schweinfurt">
          <OFFICIALS>
            <OFFICIAL officialid="23662" firstname="Andrè" gender="M" lastname="Krause" nation="GER">
              <CONTACT city="SC Schweinfurt" />
            </OFFICIAL>
            <OFFICIAL officialid="23607" firstname="Niko" gender="M" lastname="Scholz" nation="GER">
              <CONTACT city="SC Schweinfurt" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4175" nation="GER" region="02" clubid="7908" name="ASV 1860 Neumarkt" />
        <CLUB type="CLUB" code="4168" nation="GER" region="02" clubid="7962" name="ASV Cham" />
        <CLUB type="CLUB" code="4169" nation="GER" region="02" clubid="7940" name="ATS Kulmbach" />
        <CLUB type="CLUB" nation="GER" clubid="7951" name="BSV">
          <OFFICIALS>
            <OFFICIAL officialid="23560" firstname="Ingolf" gender="M" lastname="Baumbach" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23597" firstname="Julian" gender="M" lastname="Beyer" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23664" firstname="Roland" gender="M" lastname="Hanselmann" nation="GER">
              <CONTACT city="SV Dachau" />
            </OFFICIAL>
            <OFFICIAL officialid="17223" firstname="Manfred" gender="M" grade="REF" lastname="Kellner" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23581" firstname="Kerstin" gender="F" lastname="Kern" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23552" firstname="Hannes" gender="M" lastname="Kießling" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23561" firstname="Reinhard" gender="M" lastname="Kunze" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23576" firstname="Markus" gender="M" lastname="Runte" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23606" firstname="Wolfgang" gender="M" lastname="Rühl" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23551" firstname="Karsten" gender="M" lastname="Schmidt" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23594" firstname="Katja" gender="M" lastname="Scholz" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23661" firstname="Werner" gender="M" lastname="Strasser" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23660" firstname="Julia" gender="F" lastname="Strobel" nation="GER">
              <CONTACT city="SC Haßberge" />
            </OFFICIAL>
            <OFFICIAL officialid="23596" firstname="Werner" gender="M" lastname="Sturm" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23565" firstname="Roland" gender="M" lastname="Vogel" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23582" firstname="Thomas" gender="M" lastname="Weiß" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23559" firstname="Caroline" gender="M" lastname="Werner" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4224" nation="GER" region="02" clubid="7950" name="Delphin 77 Herzogenaurach">
          <OFFICIALS>
            <OFFICIAL officialid="23668" firstname="Kathrin" gender="F" lastname="Janes" nation="GER">
              <CONTACT city="Delphin Herzogenaurach" />
            </OFFICIAL>
            <OFFICIAL officialid="17215" firstname="Silke" gender="F" lastname="Janes" nation="GER">
              <CONTACT city="Delphin Herzog" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4233" nation="GER" region="02" clubid="7965" name="DJK Sportbund München" />
        <CLUB type="CLUB" code="4249" nation="GER" region="02" clubid="7959" name="FW München" />
        <CLUB type="CLUB" code="4264" nation="GER" region="02" clubid="7914" name="MTV 1862 Pfaffenhofen/Ilm" />
        <CLUB type="CLUB" code="4269" nation="GER" region="02" clubid="7954" name="Polizei SV Eichstätt" />
        <CLUB type="CLUB" code="4271" nation="GER" region="02" clubid="7892" name="Post-SV Nürnberg">
          <ATHLETES>
            <ATHLETE birthdate="2009-01-01" firstname="Helena" gender="F" lastname="Bersch" nation="GER" license="383933" athleteid="24349">
              <ENTRIES>
                <ENTRY entrytime="00:03:30.54" eventid="1183" heatid="25817" lane="2" />
                <ENTRY entrytime="00:01:49.00" eventid="1111" heatid="25850" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="1135" heatid="25894" lane="2" />
                <ENTRY entrytime="00:01:55.00" eventid="7788" heatid="25940" lane="3" />
                <ENTRY entrytime="00:00:45.00" eventid="1123" heatid="25965" lane="4" />
                <ENTRY entrytime="00:03:50.00" eventid="5661" heatid="26009" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Tobias" gender="M" lastname="Bonn" nation="GER" license="383469" athleteid="24356">
              <ENTRIES>
                <ENTRY entrytime="00:03:02.61" eventid="1177" heatid="25812" lane="4" />
                <ENTRY entrytime="00:01:36.77" eventid="1141" heatid="25885" lane="5" />
                <ENTRY entrytime="00:01:35.29" eventid="7773" heatid="25935" lane="6" />
                <ENTRY entrytime="00:01:32.37" eventid="1165" heatid="25971" lane="3" />
                <ENTRY entrytime="00:01:26.35" eventid="1189" heatid="25990" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Emilia" gender="F" lastname="Collmer" nation="GER" license="383474" athleteid="24362">
              <ENTRIES>
                <ENTRY entrytime="00:02:38.99" eventid="1183" heatid="25820" lane="3" />
                <ENTRY entrytime="00:01:37.73" eventid="1111" heatid="25851" lane="6" />
                <ENTRY entrytime="00:01:45.74" eventid="1135" heatid="25895" lane="4" />
                <ENTRY entrytime="00:01:18.85" eventid="1171" heatid="25980" lane="4" />
                <ENTRY entrytime="00:01:11.28" eventid="1195" heatid="26005" lane="3" />
                <ENTRY entrytime="00:03:02.11" eventid="5661" heatid="26011" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lukas" gender="M" lastname="Derksen" nation="GER" license="397136" athleteid="24369">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.38" eventid="5702" heatid="25828" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="1141" heatid="25883" lane="2" />
                <ENTRY entrytime="00:00:41.75" eventid="5740" heatid="25908" lane="4" />
                <ENTRY entrytime="00:00:24.46" eventid="7804" heatid="25949" lane="2" />
                <ENTRY entrytime="00:01:40.72" eventid="1189" heatid="25987" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Maxim" gender="M" lastname="Derksen" nation="GER" license="386632" athleteid="24375">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.65" eventid="5702" heatid="25832" lane="3" />
                <ENTRY entrytime="00:01:37.59" eventid="1141" heatid="25885" lane="6" />
                <ENTRY entrytime="00:00:35.71" eventid="5740" heatid="25910" lane="3" />
                <ENTRY entrytime="00:00:55.34" eventid="1117" heatid="25958" lane="1" />
                <ENTRY entrytime="00:01:22.44" eventid="1189" heatid="25991" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Tom Norman" gender="M" lastname="Dürrschmidt" nation="GER" license="386631" athleteid="24381">
              <ENTRIES>
                <ENTRY entrytime="00:02:51.27" eventid="1177" heatid="25813" lane="5" />
                <ENTRY entrytime="00:01:51.92" eventid="1141" heatid="25883" lane="6" />
                <ENTRY entrytime="00:01:44.19" eventid="7773" heatid="25934" lane="6" />
                <ENTRY entrytime="00:01:35.55" eventid="1165" heatid="25971" lane="4" />
                <ENTRY entrytime="00:01:21.48" eventid="1189" heatid="25991" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Gedion" gender="M" lastname="Efrem" nation="GER" license="392230" athleteid="24387">
              <ENTRIES>
                <ENTRY entrytime="00:03:20.66" eventid="1177" heatid="25811" lane="5" />
                <ENTRY entrytime="00:01:49.00" eventid="1103" heatid="25848" lane="5" />
                <ENTRY entrytime="00:01:45.00" eventid="7773" heatid="25933" lane="2" />
                <ENTRY entrytime="00:00:49.00" eventid="1117" heatid="25959" lane="1" />
                <ENTRY entrytime="00:01:37.00" eventid="1165" heatid="25971" lane="2" />
                <ENTRY entrytime="00:03:50.00" eventid="5655" heatid="26006" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Hasset" gender="F" lastname="Efrem" nation="GER" license="392225" athleteid="24394">
              <ENTRIES>
                <ENTRY entrytime="00:03:22.50" eventid="1183" heatid="25818" lane="1" />
                <ENTRY entrytime="00:01:57.11" eventid="1111" heatid="25849" lane="4" />
                <ENTRY entrytime="00:01:41.87" eventid="1171" heatid="25978" lane="6" />
                <ENTRY entrytime="00:01:25.67" eventid="1195" heatid="26003" lane="3" />
                <ENTRY entrytime="00:03:48.11" eventid="5661" heatid="26009" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Mathilda" gender="F" lastname="Egelkraut" nation="GER" license="399536" athleteid="24400">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="5664" heatid="25754" lane="2" />
                <ENTRY entrytime="00:00:39.00" eventid="5682" heatid="25771" lane="3" />
                <ENTRY entrytime="00:00:39.00" eventid="5690" heatid="25796" lane="5" />
                <ENTRY entrytime="00:00:48.00" eventid="5698" heatid="25804" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Nick" gender="M" lastname="Frohmeyer" nation="GER" license="394367" athleteid="24405">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.68" eventid="5702" heatid="25828" lane="5" />
                <ENTRY entrytime="00:00:53.59" eventid="5724" heatid="25859" lane="4" />
                <ENTRY entrytime="00:00:51.62" eventid="5740" heatid="25903" lane="3" />
                <ENTRY entrytime="00:01:54.97" eventid="1165" heatid="25969" lane="5" />
                <ENTRY entrytime="00:01:58.00" eventid="1189" heatid="25984" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Thomas" gender="M" lastname="Ganin" nation="GER" license="382767" athleteid="24411">
              <ENTRIES>
                <ENTRY entrytime="00:02:56.12" eventid="1177" heatid="25812" lane="3" />
                <ENTRY entrytime="00:00:33.66" eventid="5740" heatid="25911" lane="2" />
                <ENTRY entrytime="00:01:39.00" eventid="7773" heatid="25934" lane="4" />
                <ENTRY entrytime="00:00:40.89" eventid="1117" heatid="25960" lane="2" />
                <ENTRY entrytime="00:01:15.52" eventid="1189" heatid="25992" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Daniel" gender="M" lastname="Hadersbrunner" nation="GER" license="392488" athleteid="24417">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.80" eventid="5702" heatid="25827" lane="5" />
                <ENTRY entrytime="00:00:51.88" eventid="5724" heatid="25860" lane="1" />
                <ENTRY entrytime="00:00:44.49" eventid="5740" heatid="25907" lane="4" />
                <ENTRY entrytime="00:01:48.88" eventid="1165" heatid="25970" lane="5" />
                <ENTRY entrytime="00:01:40.31" eventid="1189" heatid="25987" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Marco" gender="M" lastname="Hadersbrunner" nation="GER" license="392487" athleteid="24423">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.00" eventid="5702" heatid="25829" lane="6" />
                <ENTRY entrytime="00:00:47.00" eventid="5724" heatid="25862" lane="1" />
                <ENTRY entrytime="00:00:43.38" eventid="5740" heatid="25908" lane="6" />
                <ENTRY entrytime="00:00:22.22" eventid="7804" heatid="25949" lane="3" />
                <ENTRY entrytime="00:01:45.00" eventid="1189" heatid="25986" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Simon" gender="M" lastname="Hadersbrunner" nation="GER" license="383461" athleteid="24429">
              <ENTRIES>
                <ENTRY entrytime="00:01:36.84" eventid="1103" heatid="25848" lane="3" />
                <ENTRY entrytime="00:01:41.46" eventid="1141" heatid="25884" lane="3" />
                <ENTRY entrytime="00:01:31.54" eventid="7773" heatid="25935" lane="4" />
                <ENTRY entrytime="00:00:40.13" eventid="1117" heatid="25960" lane="4" />
                <ENTRY entrytime="00:01:17.95" eventid="1189" heatid="25992" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Greta" gender="F" lastname="Haesler" nation="GER" license="383471" athleteid="24435">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.48" eventid="5712" heatid="25845" lane="3" />
                <ENTRY entrytime="00:01:47.29" eventid="1135" heatid="25895" lane="5" />
                <ENTRY entrytime="00:00:41.75" eventid="5744" heatid="25925" lane="6" />
                <ENTRY entrytime="00:01:46.16" eventid="7788" heatid="25943" lane="1" />
                <ENTRY entrytime="00:01:36.57" eventid="1195" heatid="26001" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ferdinand" gender="M" lastname="Hartmann" nation="GER" license="392484" athleteid="24441">
              <ENTRIES>
                <ENTRY entrytime="00:03:19.00" eventid="1177" heatid="25811" lane="2" />
                <ENTRY entrytime="00:00:47.35" eventid="5724" heatid="25862" lane="6" />
                <ENTRY entrytime="00:00:41.50" eventid="5740" heatid="25909" lane="6" />
                <ENTRY entrytime="00:00:19.00" eventid="7804" heatid="25950" lane="3" />
                <ENTRY entrytime="00:01:40.00" eventid="1165" heatid="25971" lane="6" />
                <ENTRY entrytime="00:01:33.44" eventid="1189" heatid="25989" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Laura" gender="F" lastname="Hartmann" nation="GER" license="383478" athleteid="24448">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.89" eventid="5712" heatid="25847" lane="5" />
                <ENTRY entrytime="00:01:47.32" eventid="1111" heatid="25850" lane="4" />
                <ENTRY entrytime="00:01:38.75" eventid="1135" heatid="25897" lane="5" />
                <ENTRY entrytime="00:01:41.05" eventid="1171" heatid="25978" lane="2" />
                <ENTRY entrytime="00:01:28.16" eventid="1195" heatid="26003" lane="4" />
                <ENTRY entrytime="00:03:23.53" eventid="5661" heatid="26011" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Leonora" gender="F" lastname="Hartmann" nation="GER" license="0" athleteid="24455">
              <ENTRIES>
                <ENTRY entrytime="00:00:35.00" eventid="5664" heatid="25754" lane="5" />
                <ENTRY entrytime="00:00:36.00" eventid="5682" heatid="25772" lane="1" />
                <ENTRY entrytime="00:00:40.00" eventid="5690" heatid="25796" lane="1" />
                <ENTRY entrytime="00:00:40.00" eventid="5698" heatid="25804" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lorenz" gender="M" lastname="Hillebrand" nation="GER" license="383463" athleteid="24460">
              <ENTRIES>
                <ENTRY entrytime="00:03:06.59" eventid="1177" heatid="25812" lane="2" />
                <ENTRY entrytime="00:01:50.24" eventid="1141" heatid="25883" lane="1" />
                <ENTRY entrytime="00:01:25.48" eventid="1165" heatid="25972" lane="5" />
                <ENTRY entrytime="00:01:23.91" eventid="1189" heatid="25990" lane="3" />
                <ENTRY entrytime="00:03:27.33" eventid="5655" heatid="26007" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="David" gender="M" lastname="Höhne" nation="GER" license="0" athleteid="24466">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.00" eventid="1053" heatid="25748" lane="2" />
                <ENTRY entrytime="00:00:41.00" eventid="5668" heatid="25759" lane="4" />
                <ENTRY entrytime="00:00:42.00" eventid="5678" heatid="25768" lane="6" />
                <ENTRY entrytime="00:00:45.00" eventid="5694" heatid="25799" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Lorenz" gender="M" lastname="Kolb" nation="GER" license="389295" athleteid="24471">
              <ENTRIES>
                <ENTRY entrytime="00:03:08.35" eventid="1177" heatid="25812" lane="5" />
                <ENTRY entrytime="00:01:49.00" eventid="1103" heatid="25848" lane="1" />
                <ENTRY entrytime="00:01:53.84" eventid="1141" heatid="25882" lane="1" />
                <ENTRY entrytime="00:01:47.65" eventid="1165" heatid="25970" lane="2" />
                <ENTRY entrytime="00:01:27.54" eventid="1189" heatid="25990" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Mathilde" gender="F" lastname="Korda" nation="GER" license="392480" athleteid="24477">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.36" eventid="5712" status="DNS" heatid="25844" lane="4" />
                <ENTRY entrytime="00:00:45.17" eventid="5728" status="DNS" heatid="25876" lane="3" />
                <ENTRY entrytime="00:00:37.39" eventid="5744" status="DNS" heatid="25927" lane="6" />
                <ENTRY entrytime="00:00:25.44" eventid="7809" status="DNS" heatid="25953" lane="3" />
                <ENTRY entrytime="00:01:24.52" eventid="1195" status="DNS" heatid="26004" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Karen" gender="F" lastname="Lothwesen" nation="GER" license="383467" athleteid="24483">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.57" eventid="5712" heatid="25847" lane="3" />
                <ENTRY entrytime="00:01:36.67" eventid="1135" heatid="25897" lane="4" />
                <ENTRY entrytime="00:00:34.44" eventid="5744" heatid="25928" lane="4" />
                <ENTRY entrytime="00:01:33.52" eventid="7788" heatid="25945" lane="2" />
                <ENTRY entrytime="00:01:24.25" eventid="1195" heatid="26004" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Elmercy" gender="F" lastname="Lulseged" nation="GER" license="0" athleteid="24489">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.00" eventid="5664" heatid="25755" lane="2" />
                <ENTRY entrytime="00:00:33.00" eventid="5682" heatid="25772" lane="2" />
                <ENTRY entrytime="00:00:34.00" eventid="5690" heatid="25796" lane="4" />
                <ENTRY entrytime="00:00:30.00" eventid="5698" heatid="25806" lane="6" />
                <ENTRY entrytime="00:00:36.00" eventid="7706" heatid="25809" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Johannes" gender="M" lastname="Lulseged" nation="GER" license="0" athleteid="24495">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.00" eventid="1053" heatid="25748" lane="5" />
                <ENTRY entrytime="00:00:48.00" eventid="5668" heatid="25759" lane="6" />
                <ENTRY entrytime="00:00:51.00" eventid="5678" heatid="25767" lane="6" />
                <ENTRY entrytime="00:00:41.00" eventid="5694" heatid="25799" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Rebekah" gender="F" lastname="Lulseged" nation="GER" license="383476" athleteid="24500">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.17" eventid="5728" heatid="25874" lane="4" />
                <ENTRY entrytime="00:00:38.77" eventid="5744" heatid="25926" lane="2" />
                <ENTRY entrytime="00:01:44.02" eventid="7788" heatid="25944" lane="6" />
                <ENTRY entrytime="00:00:50.06" eventid="1123" heatid="25963" lane="4" />
                <ENTRY entrytime="00:01:28.41" eventid="1195" heatid="26003" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Meggy" gender="F" lastname="Messel" nation="GER" license="0" athleteid="24506">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.00" eventid="5664" heatid="25755" lane="6" />
                <ENTRY entrytime="00:00:22.50" eventid="5682" heatid="25773" lane="4" />
                <ENTRY entrytime="00:00:29.00" eventid="7696" heatid="25785" lane="3" />
                <ENTRY entrytime="00:00:26.00" eventid="5698" heatid="25806" lane="4" />
                <ENTRY entrytime="00:00:28.00" eventid="7706" heatid="25809" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Michelle" gender="F" lastname="Möbus" nation="GER" license="0" athleteid="24512">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.00" eventid="5664" heatid="25755" lane="5" />
                <ENTRY entrytime="00:00:36.00" eventid="5674" heatid="25764" lane="4" />
                <ENTRY entrytime="00:00:32.00" eventid="5682" heatid="25772" lane="4" />
                <ENTRY entrytime="00:00:30.00" eventid="7696" heatid="25785" lane="4" />
                <ENTRY entrytime="00:00:36.00" eventid="5698" heatid="25805" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Sophie" gender="F" lastname="Oberndorfer" nation="GER" license="383466" athleteid="24518">
              <ENTRIES>
                <ENTRY entrytime="00:02:44.41" eventid="1183" heatid="25820" lane="2" />
                <ENTRY entrytime="00:01:26.40" eventid="1111" heatid="25851" lane="4" />
                <ENTRY entrytime="00:01:44.00" eventid="1135" heatid="25896" lane="5" />
                <ENTRY entrytime="00:01:28.00" eventid="1171" heatid="25980" lane="1" />
                <ENTRY entrytime="00:01:16.00" eventid="1195" heatid="26005" lane="4" />
                <ENTRY entrytime="00:03:14.09" eventid="5661" heatid="26011" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Sarah" gender="F" lastname="Olalowo" nation="GER" license="383462" athleteid="24525">
              <ENTRIES>
                <ENTRY entrytime="00:03:09.51" eventid="1183" heatid="25818" lane="3" />
                <ENTRY entrytime="00:00:42.61" eventid="5712" heatid="25847" lane="4" />
                <ENTRY entrytime="00:01:30.53" eventid="1135" heatid="25897" lane="3" />
                <ENTRY entrytime="00:01:40.00" eventid="7788" heatid="25944" lane="2" />
                <ENTRY entrytime="00:01:37.21" eventid="1171" heatid="25979" lane="6" />
                <ENTRY entrytime="00:01:24.72" eventid="1195" heatid="26004" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Alexander" gender="M" lastname="Primorac" nation="GER" license="392226" athleteid="24532">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.97" eventid="5702" heatid="25831" lane="3" />
                <ENTRY entrytime="00:01:48.63" eventid="1141" heatid="25884" lane="6" />
                <ENTRY entrytime="00:01:40.00" eventid="7773" heatid="25934" lane="5" />
                <ENTRY entrytime="00:01:45.00" eventid="1165" heatid="25970" lane="4" />
                <ENTRY entrytime="00:01:25.62" eventid="1189" heatid="25990" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Carla" gender="F" lastname="Primorac" nation="GER" license="392227" athleteid="24538">
              <ENTRIES>
                <ENTRY entrytime="00:03:13.86" eventid="1183" heatid="25818" lane="4" />
                <ENTRY entrytime="00:01:57.71" eventid="1135" heatid="25893" lane="6" />
                <ENTRY entrytime="00:00:46.27" eventid="1123" heatid="25965" lane="1" />
                <ENTRY entrytime="00:01:41.72" eventid="1171" heatid="25978" lane="1" />
                <ENTRY entrytime="00:01:30.98" eventid="1195" heatid="26002" lane="4" />
                <ENTRY entrytime="00:03:35.46" eventid="5661" heatid="26010" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Elijas" gender="M" lastname="Rau" nation="GER" license="397135" athleteid="24545">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.69" eventid="5702" heatid="25826" lane="2" />
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25881" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5740" heatid="25904" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Nick" gender="M" lastname="Rein" nation="GER" license="416115" athleteid="24549">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5702" heatid="25825" lane="6" />
                <ENTRY entrytime="00:01:04.00" eventid="5724" heatid="25855" lane="5" />
                <ENTRY entrytime="00:00:50.98" eventid="5740" heatid="25904" lane="6" />
                <ENTRY entrytime="00:00:35.00" eventid="7804" heatid="25947" lane="5" />
                <ENTRY entrytime="00:01:58.07" eventid="1189" heatid="25984" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Clara" gender="F" lastname="Seibold" nation="GER" license="0" athleteid="24555">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.00" eventid="5664" heatid="25754" lane="6" />
                <ENTRY entrytime="00:00:39.00" eventid="5682" heatid="25771" lane="4" />
                <ENTRY entrytime="00:00:41.00" eventid="5690" heatid="25796" lane="6" />
                <ENTRY entrytime="00:00:43.00" eventid="5698" heatid="25804" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Henry" gender="M" lastname="Shi" nation="GER" license="393061" athleteid="24560">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.72" eventid="5702" heatid="25830" lane="3" />
                <ENTRY entrytime="00:00:48.42" eventid="5724" heatid="25861" lane="3" />
                <ENTRY entrytime="00:01:53.53" eventid="1141" heatid="25882" lane="2" />
                <ENTRY entrytime="00:00:22.04" eventid="7804" heatid="25950" lane="6" />
                <ENTRY entrytime="00:01:31.98" eventid="1189" heatid="25989" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Nea" gender="F" lastname="Stöckel" nation="GER" license="382760" athleteid="24566">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.92" eventid="1183" heatid="25820" lane="1" />
                <ENTRY entrytime="00:01:29.00" eventid="1111" heatid="25851" lane="5" />
                <ENTRY entrytime="00:01:40.00" eventid="1135" heatid="25897" lane="6" />
                <ENTRY entrytime="00:00:39.08" eventid="1123" heatid="25966" lane="4" />
                <ENTRY entrytime="00:01:16.43" eventid="1195" heatid="26005" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Maximilian" gender="M" lastname="Tatár" nation="GER" license="412059" athleteid="24572">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5702" heatid="25824" lane="3" />
                <ENTRY entrytime="00:01:05.00" eventid="5724" heatid="25855" lane="6" />
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25881" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5740" heatid="25901" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lukas" gender="M" lastname="Westphal" nation="GER" license="412060" athleteid="24577">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.29" eventid="5724" status="DNS" heatid="25859" lane="6" />
                <ENTRY entrytime="00:00:46.99" eventid="5740" heatid="25906" lane="5" />
                <ENTRY entrytime="00:00:33.00" eventid="7804" heatid="25947" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="1165" heatid="25970" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Arnold" gender="M" lastname="Zinoviev" nation="GER" license="412058" athleteid="24582">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.00" eventid="5702" heatid="25832" lane="5" />
                <ENTRY entrytime="00:01:50.00" eventid="1141" heatid="25883" lane="3" />
                <ENTRY entrytime="00:00:45.00" eventid="5740" heatid="25907" lane="5" />
                <ENTRY entrytime="00:00:20.00" eventid="7804" heatid="25950" lane="4" />
                <ENTRY entrytime="00:00:52.00" eventid="1117" heatid="25958" lane="5" />
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25986" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="8" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:02:27.69" eventid="23774" heatid="25946" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="24460" number="1" />
                    <RELAYPOSITION athleteid="24483" number="2" />
                    <RELAYPOSITION athleteid="24566" number="3" />
                    <RELAYPOSITION athleteid="24411" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="23767" firstname="Doris" gender="F" lastname="Colmer" nation="GER">
              <CONTACT city="Post SV Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="17212" firstname="Nicole" gender="F" lastname="Hadersbrunner" nation="GER">
              <CONTACT city="Post-SV Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="17185" firstname="Liane" gender="F" lastname="Hindelang" nation="GER">
              <CONTACT city="Post SV Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="26098" firstname="Christian" gender="M" lastname="Korda" nation="GER">
              <CONTACT city="Post-SV Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="23655" firstname="Steffi" gender="M" lastname="Korda" nation="GER">
              <CONTACT city="Post SV Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="23667" firstname="Marlies" gender="F" lastname="Lifka" nation="GER">
              <CONTACT city="Post SV Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="17208" firstname="Alfred" gender="M" lastname="Seelmann" nation="GER">
              <CONTACT city="BSV" />
            </OFFICIAL>
            <OFFICIAL officialid="23665" firstname="Roswitha" gender="M" lastname="Seelmann" nation="GER">
              <CONTACT city="Post SV Nürnbaerg" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4300" nation="GER" region="02" clubid="25172" name="Sb Bayern 07">
          <ATHLETES>
            <ATHLETE birthdate="2009-01-01" firstname="Karla" gender="F" lastname="Gottwald" nation="GER" license="407071" athleteid="25173">
              <ENTRIES>
                <ENTRY entrytime="00:03:55.60" eventid="1183" heatid="25816" lane="4" />
                <ENTRY entrytime="00:01:04.10" eventid="5728" heatid="25869" lane="6" />
                <ENTRY entrytime="00:01:05.68" eventid="5744" heatid="25915" lane="6" />
                <ENTRY entrytime="00:01:30.01" eventid="1123" heatid="25961" lane="3" />
                <ENTRY entrytime="00:02:14.67" eventid="1171" heatid="25974" lane="2" />
                <ENTRY entrytime="00:02:15.15" eventid="1195" heatid="25994" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Leni" gender="F" lastname="Kreß" nation="GER" license="420601" athleteid="25180">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.32" eventid="5712" heatid="25842" lane="4" />
                <ENTRY entrytime="00:02:02.78" eventid="1135" heatid="25891" lane="5" />
                <ENTRY entrytime="00:00:56.32" eventid="5744" status="DNS" heatid="25918" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Carla-Sophie" gender="F" lastname="Lindner" nation="GER" license="407066" athleteid="25184">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.66" eventid="5712" status="DNS" heatid="25838" lane="5" />
                <ENTRY entrytime="00:01:10.20" eventid="5728" status="DNS" heatid="25866" lane="1" />
                <ENTRY entrytime="00:02:17.22" eventid="1135" status="DNS" heatid="25890" lane="5" />
                <ENTRY entrytime="00:01:10.02" eventid="5744" status="DNS" heatid="25914" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Amelie" gender="F" lastname="Maußner" nation="GER" license="420602" athleteid="25189">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25834" lane="1" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25887" lane="1" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25912" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Adrian" gender="M" lastname="Neumann" nation="GER" license="420606" athleteid="25193">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5702" heatid="25821" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Oleg" gender="M" lastname="Orazmagomedor" nation="GER" license="0" athleteid="25195">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.08" eventid="1053" status="DNS" heatid="25745" lane="4" />
                <ENTRY entrytime="NT" eventid="5686" status="DNS" heatid="25788" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ida" gender="F" lastname="Pfeuffer" nation="GER" license="407068" athleteid="25199">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.20" eventid="5728" heatid="25866" lane="6" />
                <ENTRY entrytime="00:01:07.02" eventid="5744" heatid="25914" lane="3" />
                <ENTRY entrytime="00:02:37.33" eventid="7788" heatid="25937" lane="4" />
                <ENTRY entrytime="00:01:10.14" eventid="7809" heatid="25952" lane="6" />
                <ENTRY entrytime="00:02:15.00" eventid="1171" heatid="25974" lane="5" />
                <ENTRY entrytime="00:02:13.00" eventid="1195" heatid="25995" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Lisa" gender="F" lastname="Richter" nation="GER" license="0" athleteid="25206">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.67" eventid="5664" heatid="25752" lane="6" />
                <ENTRY entrytime="00:00:55.67" eventid="5682" heatid="25770" lane="3" />
                <ENTRY entrytime="00:01:23.39" eventid="7696" heatid="25783" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Vivien-Sarah" gender="F" lastname="Richter" nation="GER" license="407525" athleteid="25210">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.20" eventid="5712" heatid="25838" lane="1" />
                <ENTRY entrytime="00:01:03.20" eventid="5728" heatid="25869" lane="2" />
                <ENTRY entrytime="00:02:18.67" eventid="1135" heatid="25890" lane="6" />
                <ENTRY entrytime="00:00:58.18" eventid="5744" heatid="25917" lane="3" />
                <ENTRY entrytime="00:02:13.22" eventid="1171" heatid="25974" lane="4" />
                <ENTRY entrytime="00:02:03.36" eventid="1195" heatid="25996" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Felix" gender="M" lastname="Schäfer" nation="GER" license="0" athleteid="25217">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.17" eventid="1053" heatid="25746" lane="4" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25775" lane="6" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25789" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Jakob" gender="M" lastname="Schäfer" nation="GER" license="420605" athleteid="25221">
              <ENTRIES>
                <ENTRY entrytime="00:01:19.41" eventid="5702" heatid="25822" lane="2" />
                <ENTRY entrytime="00:02:45.41" eventid="1141" heatid="25878" lane="3" />
                <ENTRY entrytime="00:01:15.67" eventid="5740" heatid="25900" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Nils" gender="M" lastname="Wunderlich" nation="GER" license="420599" athleteid="25225">
              <ENTRIES>
                <ENTRY entrytime="00:03:40.20" eventid="1177" heatid="25810" lane="4" />
                <ENTRY entrytime="00:01:03.03" eventid="5724" heatid="25855" lane="2" />
                <ENTRY entrytime="00:00:46.20" eventid="5740" heatid="25906" lane="4" />
                <ENTRY entrytime="00:02:15.20" eventid="7773" heatid="25930" lane="3" />
                <ENTRY entrytime="00:02:10.10" eventid="1165" heatid="25968" lane="1" />
                <ENTRY entrytime="00:01:55.66" eventid="1189" heatid="25984" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Tim" gender="M" lastname="Wunderlich" nation="GER" license="420600" athleteid="25232">
              <ENTRIES>
                <ENTRY entrytime="00:01:20.00" eventid="5702" status="DNS" heatid="25822" lane="5" />
                <ENTRY entrytime="00:01:20.00" eventid="5724" status="DNS" heatid="25854" lane="1" />
                <ENTRY entrytime="00:02:45.00" eventid="1141" status="DNS" heatid="25879" lane="6" />
                <ENTRY entrytime="00:01:16.00" eventid="5740" status="DNS" heatid="25900" lane="1" />
                <ENTRY entrytime="00:02:40.80" eventid="1165" status="DNS" heatid="25967" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Charlotte" gender="F" lastname="Zimmermann" nation="GER" license="420604" athleteid="25238">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.20" eventid="5712" status="DNS" heatid="25838" lane="6" />
                <ENTRY entrytime="00:01:04.54" eventid="5728" status="DNS" heatid="25868" lane="3" />
                <ENTRY entrytime="00:02:20.20" eventid="1135" status="DNS" heatid="25889" lane="5" />
                <ENTRY entrytime="00:01:10.70" eventid="5744" status="DNS" heatid="25914" lane="1" />
                <ENTRY entrytime="00:02:16.20" eventid="1171" status="DNS" heatid="25973" lane="3" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4280" nation="GER" region="02" clubid="7972" name="SB Delphin 03 Augsburg" />
        <CLUB type="CLUB" code="4290" nation="GER" region="02" clubid="7919" name="SC 53 Landshut" />
        <CLUB type="CLUB" code="4286" nation="GER" region="02" clubid="7953" name="SC Delphin Ingolstadt" />
        <CLUB type="CLUB" code="4292" nation="GER" region="02" clubid="7974" name="SC Prinz Eugen München">
          <OFFICIALS>
            <OFFICIAL officialid="23677" firstname="Uli" gender="M" lastname="Fischer" nation="GER">
              <CONTACT city="SC Prinz Eugen M" />
            </OFFICIAL>
            <OFFICIAL officialid="23580" firstname="Uli" gender="M" lastname="Fischer" nation="GER">
              <CONTACT city="SC PE München" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="6524" nation="GER" region="02" clubid="7970" name="SC Regensburg">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="Albert" gender="M" lastname="Ackbarow" nation="GER" license="000000" athleteid="24590">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.70" eventid="5668" heatid="25760" lane="3" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25766" lane="5" />
                <ENTRY entrytime="00:00:33.30" eventid="7691" heatid="25779" lane="3" />
                <ENTRY entrytime="00:00:28.56" eventid="5694" heatid="25801" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Louis" gender="M" lastname="Bär" nation="GER" license="000000" athleteid="24595">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.89" eventid="1053" heatid="25748" lane="4" />
                <ENTRY entrytime="00:00:46.60" eventid="5668" heatid="25759" lane="1" />
                <ENTRY entrytime="00:00:34.80" eventid="7691" heatid="25779" lane="2" />
                <ENTRY entrytime="00:00:35.50" eventid="5686" heatid="25791" lane="4" />
                <ENTRY entrytime="00:00:36.11" eventid="5694" heatid="25800" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Jannik" gender="M" lastname="De Swart" nation="GER" license="000000" athleteid="24601">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25744" lane="2" />
                <ENTRY entrytime="NT" eventid="5668" heatid="25757" lane="5" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25774" lane="1" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25789" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Fabian" gender="M" lastname="Frizler" nation="GER" license="000000" athleteid="24606">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25757" lane="3" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25775" lane="2" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25787" lane="3" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25798" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Felix" gender="M" lastname="Gallner" nation="GER" license="000000" athleteid="24611">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25757" lane="2" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25774" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Helena" gender="F" lastname="Glas" nation="GER" license="000000" athleteid="24614">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25750" lane="3" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25761" lane="4" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25780" lane="2" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25792" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Leni" gender="F" lastname="Haubner" nation="GER" license="000000" athleteid="24619">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25750" lane="5" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25762" lane="1" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25781" lane="5" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25794" lane="1" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25802" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lilli" gender="F" lastname="Heindl" nation="GER" license="000000" athleteid="24625">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25751" lane="1" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25762" lane="5" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25781" lane="2" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25794" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Bruno" gender="M" lastname="Hubert" nation="GER" license="000000" athleteid="24630">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25757" lane="4" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25774" lane="4" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25787" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Johanna" gender="F" lastname="Kapfenberger" nation="GER" license="000000" athleteid="24634">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.60" eventid="5674" heatid="25764" lane="1" />
                <ENTRY entrytime="00:00:41.30" eventid="7696" heatid="25784" lane="3" />
                <ENTRY entrytime="00:00:55.30" eventid="5690" heatid="25795" lane="1" />
                <ENTRY entrytime="00:00:39.20" eventid="5698" heatid="25805" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Roman" gender="M" lastname="Kuldyaev" nation="GER" license="000000" athleteid="24645">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25756" lane="4" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25774" lane="2" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25797" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Felix" gender="M" lastname="Kübler" nation="GER" license="000000" athleteid="24639">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.30" eventid="5668" heatid="25760" lane="5" />
                <ENTRY entrytime="00:00:35.17" eventid="5678" heatid="25768" lane="4" />
                <ENTRY entrytime="00:00:36.50" eventid="7691" heatid="25779" lane="1" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25788" lane="5" />
                <ENTRY entrytime="00:00:31.80" eventid="5694" heatid="25801" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="David" gender="M" lastname="Metreveli" nation="GER" license="000000" athleteid="24649">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25757" lane="1" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25774" lane="6" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25798" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Raúl" gender="M" lastname="Muñoz" nation="GER" license="000000" athleteid="24653">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5668" heatid="25757" lane="6" />
                <ENTRY entrytime="NT" eventid="7691" status="DNS" heatid="25776" lane="4" />
                <ENTRY entrytime="NT" eventid="5686" status="DNS" heatid="25786" lane="2" />
                <ENTRY entrytime="NT" eventid="5694" status="DNS" heatid="25797" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Maya Zoe" gender="F" lastname="Orth" nation="GER" license="000000" athleteid="24658">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.95" eventid="5664" heatid="25753" lane="3" />
                <ENTRY entrytime="00:00:42.90" eventid="5674" heatid="25764" lane="6" />
                <ENTRY entrytime="00:00:46.80" eventid="5682" heatid="25771" lane="1" />
                <ENTRY entrytime="00:00:49.70" eventid="5690" heatid="25795" lane="3" />
                <ENTRY entrytime="00:00:37.24" eventid="5698" heatid="25805" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Mia" gender="F" lastname="Pauly" nation="GER" license="000000" athleteid="24664">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25750" lane="2" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25761" lane="2" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25782" lane="1" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25793" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Felix" gender="M" lastname="Ramsauer" nation="GER" license="000000" athleteid="24669">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.30" eventid="5668" heatid="25758" lane="4" />
                <ENTRY entrytime="00:00:43.50" eventid="7691" heatid="25778" lane="5" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25787" lane="4" />
                <ENTRY entrytime="00:00:52.08" eventid="5694" heatid="25799" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Leon" gender="M" lastname="Rauscher" nation="GER" license="000000" athleteid="24674">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.70" eventid="5668" heatid="25758" lane="3" />
                <ENTRY entrytime="00:00:44.30" eventid="7691" heatid="25778" lane="1" />
                <ENTRY entrytime="00:01:15.00" eventid="5686" heatid="25789" lane="4" />
                <ENTRY entrytime="00:00:49.04" eventid="5694" heatid="25799" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Marc" gender="M" lastname="Rohrmüller" nation="GER" license="000000" athleteid="24679">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.90" eventid="5668" heatid="25759" lane="3" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25766" lane="1" />
                <ENTRY entrytime="00:00:33.90" eventid="7691" heatid="25779" lane="4" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25787" lane="6" />
                <ENTRY entrytime="00:00:33.54" eventid="5694" heatid="25800" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Sebastian" gender="M" lastname="Schmid" nation="GER" license="000000" athleteid="24685">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.80" eventid="5668" heatid="25760" lane="6" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25765" lane="2" />
                <ENTRY entrytime="00:00:41.20" eventid="7691" heatid="25778" lane="3" />
                <ENTRY entrytime="00:00:45.40" eventid="5686" heatid="25791" lane="6" />
                <ENTRY entrytime="00:00:37.80" eventid="5694" heatid="25800" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Maximilian" gender="M" lastname="Siege" nation="GER" license="000000" athleteid="24691">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25745" lane="1" />
                <ENTRY entrytime="NT" eventid="5668" heatid="25756" lane="3" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25775" lane="1" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25788" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lina" gender="F" lastname="Sinkel" nation="GER" license="000000" athleteid="24696">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5674" heatid="25762" lane="4" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25780" lane="3" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25794" lane="3" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25802" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Özüm" gender="F" lastname="Yigit" nation="GER" license="000000" athleteid="24701">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5674" heatid="25762" lane="2" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25783" lane="6" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25802" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="26064" firstname="Manfred" gender="M" lastname="Kammerer" nation="GER">
              <CONTACT city="SC Regensburg" />
            </OFFICIAL>
            <OFFICIAL officialid="26068" firstname="Katja" gender="F" lastname="Kapfenberger" nation="GER">
              <CONTACT city="SC Regensburg" />
            </OFFICIAL>
            <OFFICIAL officialid="26047" firstname="Antonia" gender="F" lastname="Kirchhoff" nation="GER">
              <CONTACT city="SC Regensburg" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4383" nation="GER" region="02" clubid="7883" name="SC Uttenreuth">
          <ATHLETES>
            <ATHLETE birthdate="2009-01-01" firstname="Mariella" gender="F" lastname="Braun" nation="GER" license="414988" athleteid="25416">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5712" heatid="25839" lane="1" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25867" lane="2" />
                <ENTRY entrytime="00:01:05.00" eventid="5744" heatid="25915" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Michael" gender="M" lastname="Dittrich" nation="GER" license="000000" athleteid="25420">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.00" eventid="5678" heatid="25767" lane="3" />
                <ENTRY entrytime="00:00:55.00" eventid="7691" heatid="25777" lane="2" />
                <ENTRY entrytime="00:00:50.00" eventid="5686" heatid="25790" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Finnja" gender="F" lastname="Friederich" nation="GER" license="000000" athleteid="25424">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.00" eventid="5712" heatid="25840" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5728" heatid="25870" lane="5" />
                <ENTRY entrytime="00:01:58.00" eventid="1135" heatid="25892" lane="4" />
                <ENTRY entrytime="00:00:58.00" eventid="5744" heatid="25918" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Paul" gender="M" lastname="Glanz" nation="GER" license="000000" athleteid="25429">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.00" eventid="1053" heatid="25747" lane="3" />
                <ENTRY entrytime="00:00:38.00" eventid="5678" heatid="25768" lane="5" />
                <ENTRY entrytime="00:00:47.00" eventid="5686" heatid="25790" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Leefke" gender="F" lastname="Heyken" nation="GER" license="414984" athleteid="25433">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25836" lane="1" />
                <ENTRY entrytime="00:01:20.00" eventid="5728" heatid="25865" lane="2" />
                <ENTRY entrytime="00:01:10.00" eventid="5744" heatid="25914" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Maret" gender="F" lastname="Koller" nation="GER" license="000000" athleteid="25437">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="5664" status="DNS" heatid="25753" lane="2" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" status="DNS" heatid="25784" lane="1" />
                <ENTRY entrytime="00:00:52.00" eventid="5690" status="DNS" heatid="25795" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Alina" gender="F" lastname="Sahinbegovic" nation="GER" license="000000" athleteid="25441">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="5664" status="DNS" heatid="25753" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" status="DNS" heatid="25783" lane="3" />
                <ENTRY entrytime="00:00:52.00" eventid="5690" status="DNS" heatid="25795" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Caroline" gender="F" lastname="Wendt" nation="GER" license="000000" athleteid="25445">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="5712" heatid="25843" lane="5" />
                <ENTRY entrytime="00:00:58.00" eventid="5728" heatid="25870" lane="3" />
                <ENTRY entrytime="00:01:56.00" eventid="1135" heatid="25893" lane="1" />
                <ENTRY entrytime="00:00:58.00" eventid="5744" heatid="25918" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Sebastian" gender="M" lastname="Wendt" nation="GER" license="000000" athleteid="25450">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.00" eventid="5702" heatid="25826" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5724" heatid="25856" lane="1" />
                <ENTRY entrytime="00:01:58.00" eventid="1141" heatid="25881" lane="2" />
                <ENTRY entrytime="00:00:58.00" eventid="5740" heatid="25902" lane="2" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="17200" firstname="Anna" gender="F" lastname="Dittrich" nation="GER" />
            <OFFICIAL officialid="17199" firstname="Nils" gender="M" lastname="Dittrich" nation="GER" />
            <OFFICIAL officialid="26060" firstname="Annika" gender="F" lastname="Wallerer" nation="GER">
              <CONTACT city="SC Uttenreuth" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4296" nation="GER" region="02" clubid="7912" name="SC Wfr. München" />
        <CLUB type="CLUB" code="4298" nation="GER" region="02" clubid="7907" name="SC Zwiesel" />
        <CLUB type="CLUB" code="6777" nation="GER" region="02" clubid="23892" name="Schwimmclub Schwandorf">
          <ATHLETES>
            <ATHLETE birthdate="2012-01-01" firstname="Luca" gender="M" lastname="Daucher" nation="GER" license="404783" athleteid="23893">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.50" eventid="1053" heatid="25747" lane="6" />
                <ENTRY entrytime="00:00:44.58" eventid="5678" heatid="25767" lane="2" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25776" lane="5" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25787" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Carlotta" gender="F" lastname="Fleischmann" nation="GER" license="374674" athleteid="23898">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.64" eventid="5712" heatid="25839" lane="3" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25886" lane="3" />
                <ENTRY entrytime="00:00:59.81" eventid="5744" heatid="25917" lane="2" />
                <ENTRY entrytime="NT" eventid="7788" heatid="25936" lane="3" />
                <ENTRY entrytime="00:00:33.83" eventid="7809" heatid="25952" lane="2" />
                <ENTRY entrytime="00:02:01.38" eventid="1195" heatid="25996" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Lucie" gender="F" lastname="Gebele" nation="GER" license="405006" athleteid="23912">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.89" eventid="5664" heatid="25752" lane="3" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25761" lane="3" />
                <ENTRY entrytime="00:00:41.11" eventid="5682" heatid="25771" lane="2" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25782" lane="3" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25794" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lina-Marie" gender="F" lastname="Grünauer" nation="GER" license="420366" athleteid="23918">
              <ENTRIES>
                <ENTRY entrytime="00:05:24.93" eventid="1183" heatid="25815" lane="5" />
                <ENTRY entrytime="00:01:05.13" eventid="5712" heatid="25837" lane="5" />
                <ENTRY entrytime="NT" eventid="1135" status="DNS" heatid="25888" lane="6" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25912" lane="5" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25951" lane="5" />
                <ENTRY entrytime="NT" eventid="1171" heatid="25973" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Helena" gender="F" lastname="Gäntzle" nation="GER" license="405005" athleteid="23905">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25833" lane="3" />
                <ENTRY entrytime="NT" eventid="5728" heatid="25864" lane="2" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25887" lane="5" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25912" lane="4" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25951" lane="4" />
                <ENTRY entrytime="NT" eventid="1195" heatid="25993" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Hannah" gender="F" lastname="Hecht" nation="GER" license="374659" athleteid="23925">
              <ENTRIES>
                <ENTRY entrytime="00:03:41.41" eventid="1183" heatid="25817" lane="5" />
                <ENTRY entrytime="00:00:51.04" eventid="5712" status="DNS" heatid="25844" lane="3" />
                <ENTRY entrytime="00:01:53.10" eventid="1135" status="DNS" heatid="25893" lane="3" />
                <ENTRY entrytime="NT" eventid="7788" status="DNS" heatid="25937" lane="5" />
                <ENTRY entrytime="00:01:04.37" eventid="1123" status="DNS" heatid="25962" lane="1" />
                <ENTRY entrytime="00:01:40.29" eventid="1195" status="DNS" heatid="26001" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Andreas" gender="M" lastname="Hiltl" nation="GER" license="371456" athleteid="23932">
              <ENTRIES>
                <ENTRY entrytime="00:05:01.89" eventid="1177" heatid="25810" lane="1" />
                <ENTRY entrytime="NT" eventid="1141" heatid="25878" lane="4" />
                <ENTRY entrytime="00:00:48.53" eventid="5740" heatid="25904" lane="3" />
                <ENTRY entrytime="00:02:50.44" eventid="7773" heatid="25930" lane="4" />
                <ENTRY entrytime="00:00:30.96" eventid="7804" heatid="25947" lane="3" />
                <ENTRY entrytime="00:01:59.14" eventid="1189" heatid="25984" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emma" gender="F" lastname="Knerer" nation="GER" license="374660" athleteid="23939">
              <ENTRIES>
                <ENTRY entrytime="00:03:59.89" eventid="1183" heatid="25816" lane="1" />
                <ENTRY entrytime="00:02:28.96" eventid="1135" heatid="25888" lane="3" />
                <ENTRY entrytime="00:00:50.31" eventid="5744" heatid="25920" lane="4" />
                <ENTRY entrytime="00:02:20.85" eventid="7788" heatid="25938" lane="4" />
                <ENTRY entrytime="NT" eventid="1123" heatid="25961" lane="2" />
                <ENTRY entrytime="00:01:55.59" eventid="1195" heatid="25998" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lena" gender="F" lastname="Knerer" nation="GER" license="404785" athleteid="23946">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.78" eventid="5664" heatid="25752" lane="4" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25780" lane="4" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25794" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emma" gender="F" lastname="Köhn" nation="GER" license="418818" athleteid="23950">
              <ENTRIES>
                <ENTRY entrytime="00:05:02.09" eventid="1183" heatid="25815" lane="2" />
                <ENTRY entrytime="NT" eventid="5728" heatid="25865" lane="6" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25912" lane="3" />
                <ENTRY entrytime="NT" eventid="7788" heatid="25936" lane="4" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25951" lane="3" />
                <ENTRY entrytime="00:02:20.24" eventid="1195" heatid="25994" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Heike" gender="F" lastname="Lanzl" nation="GER" license="390305" athleteid="23957">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.44" eventid="5712" heatid="25841" lane="1" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25887" lane="3" />
                <ENTRY entrytime="00:00:51.90" eventid="5744" heatid="25920" lane="1" />
                <ENTRY entrytime="00:02:27.15" eventid="7788" heatid="25938" lane="1" />
                <ENTRY entrytime="NT" eventid="1123" heatid="25961" lane="5" />
                <ENTRY entrytime="00:02:09.33" eventid="1195" heatid="25995" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Abby" gender="F" lastname="Lukas" nation="GER" license="374673" athleteid="23964">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.06" eventid="5712" heatid="25837" lane="2" />
                <ENTRY entrytime="00:01:03.34" eventid="5728" heatid="25869" lane="1" />
                <ENTRY entrytime="00:01:02.64" eventid="5744" heatid="25916" lane="1" />
                <ENTRY entrytime="00:02:35.30" eventid="7788" heatid="25937" lane="3" />
                <ENTRY entrytime="NT" eventid="1123" heatid="25961" lane="4" />
                <ENTRY entrytime="00:01:57.18" eventid="1195" heatid="25997" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Max" gender="M" lastname="Maderer" nation="GER" license="374755" athleteid="23971">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.86" eventid="5702" heatid="25825" lane="3" />
                <ENTRY entrytime="00:01:00.87" eventid="5724" heatid="25856" lane="6" />
                <ENTRY entrytime="00:02:20.11" eventid="1141" heatid="25879" lane="2" />
                <ENTRY entrytime="00:01:02.35" eventid="5740" heatid="25901" lane="2" />
                <ENTRY entrytime="NT" eventid="1165" heatid="25967" lane="4" />
                <ENTRY entrytime="00:02:38.43" eventid="1189" heatid="25981" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Aleksei" gender="M" lastname="Malikoski" nation="GER" license="390306" athleteid="23978">
              <ENTRIES>
                <ENTRY entrytime="00:03:34.02" eventid="1177" status="DNS" heatid="25810" lane="3" />
                <ENTRY entrytime="00:00:59.83" eventid="5724" status="DNS" heatid="25856" lane="2" />
                <ENTRY entrytime="00:00:47.62" eventid="5740" status="DNS" heatid="25906" lane="6" />
                <ENTRY entrytime="NT" eventid="7773" status="DNS" heatid="25929" lane="3" />
                <ENTRY entrytime="00:01:04.38" eventid="1117" status="DNS" heatid="25957" lane="1" />
                <ENTRY entrytime="00:01:36.83" eventid="1189" status="DNS" heatid="25988" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Eva" gender="F" lastname="Matthes" nation="GER" license="000000" athleteid="23985">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.04" eventid="5664" heatid="25752" lane="5" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25782" lane="4" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25793" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Ida" gender="F" lastname="Matthes" nation="GER" license="416783" athleteid="23989">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.71" eventid="5712" heatid="25835" lane="5" />
                <ENTRY entrytime="NT" eventid="5728" heatid="25864" lane="5" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25886" lane="2" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25913" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Hanna" gender="F" lastname="Rieder" nation="GER" license="390308" athleteid="23995">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.19" eventid="5712" heatid="25837" lane="1" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25888" lane="1" />
                <ENTRY entrytime="00:01:07.79" eventid="5744" heatid="25914" lane="4" />
                <ENTRY entrytime="00:02:44.76" eventid="7788" heatid="25937" lane="2" />
                <ENTRY entrytime="NT" eventid="1123" heatid="25961" lane="1" />
                <ENTRY entrytime="00:02:10.62" eventid="1195" heatid="25995" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="David" gender="M" lastname="Schlundt" nation="GER" license="390309" athleteid="24002">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.46" eventid="1053" heatid="25748" lane="6" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25766" lane="2" />
                <ENTRY entrytime="NT" eventid="7691" status="DNS" heatid="25774" lane="5" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25787" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leonie" gender="F" lastname="Seger" nation="GER" license="390311" athleteid="24007">
              <ENTRIES>
                <ENTRY entrytime="00:03:53.14" eventid="1183" heatid="25816" lane="3" />
                <ENTRY entrytime="00:00:55.01" eventid="5728" heatid="25872" lane="1" />
                <ENTRY entrytime="00:00:51.28" eventid="5744" heatid="25920" lane="5" />
                <ENTRY entrytime="00:02:23.25" eventid="7788" heatid="25938" lane="5" />
                <ENTRY entrytime="00:00:24.30" eventid="7809" heatid="25954" lane="5" />
                <ENTRY entrytime="00:01:51.95" eventid="1195" heatid="25998" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Zoe" gender="F" lastname="Seger" nation="GER" license="390312" athleteid="24014">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.31" eventid="5664" heatid="25755" lane="1" />
                <ENTRY entrytime="00:00:21.34" eventid="5682" heatid="25773" lane="3" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25781" lane="1" />
                <ENTRY entrytime="00:00:27.18" eventid="5698" heatid="25806" lane="5" />
                <ENTRY entrytime="NT" eventid="7706" heatid="25808" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Anton" gender="M" lastname="Stiegler" nation="GER" license="000000" athleteid="24020">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.51" eventid="1053" heatid="25746" lane="3" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25775" lane="3" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25786" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lara" gender="F" lastname="Wachtel" nation="GER" license="404786" athleteid="24024">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.75" eventid="5664" heatid="25753" lane="4" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25762" lane="6" />
                <ENTRY entrytime="00:00:37.65" eventid="5682" heatid="25772" lane="6" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25781" lane="4" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25794" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lea" gender="F" lastname="Wachtel" nation="GER" license="374672" athleteid="24030">
              <ENTRIES>
                <ENTRY entrytime="00:04:20.49" eventid="1183" heatid="25815" lane="3" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25888" lane="2" />
                <ENTRY entrytime="00:00:47.97" eventid="5744" heatid="25922" lane="1" />
                <ENTRY entrytime="00:02:22.04" eventid="7788" heatid="25938" lane="2" />
                <ENTRY entrytime="00:00:27.99" eventid="7809" heatid="25953" lane="6" />
                <ENTRY entrytime="00:01:53.06" eventid="1195" heatid="25998" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Emil" gender="M" lastname="Wiederer" nation="GER" license="404787" athleteid="24037">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.50" eventid="1053" heatid="25746" lane="2" />
                <ENTRY entrytime="00:00:44.58" eventid="5678" heatid="25767" lane="5" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25776" lane="2" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25788" lane="4" />
                <ENTRY entrytime="NT" eventid="7701" heatid="25807" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Pauline" gender="F" lastname="Wiederer" nation="GER" license="390242" athleteid="24043">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.95" eventid="5712" heatid="25838" lane="3" />
                <ENTRY entrytime="00:02:17.44" eventid="1135" heatid="25890" lane="1" />
                <ENTRY entrytime="00:02:32.38" eventid="7788" heatid="25938" lane="6" />
                <ENTRY entrytime="00:00:26.40" eventid="7809" heatid="25953" lane="1" />
                <ENTRY entrytime="00:02:11.24" eventid="1171" heatid="25975" lane="6" />
                <ENTRY entrytime="00:02:11.56" eventid="1195" heatid="25995" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Emma" gender="F" lastname="Zausinger" nation="GER" license="390314" athleteid="24050">
              <ENTRIES>
                <ENTRY entrytime="00:04:39.00" eventid="1183" heatid="25815" lane="4" />
                <ENTRY entrytime="00:01:11.74" eventid="5712" heatid="25835" lane="4" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25886" lane="4" />
                <ENTRY entrytime="NT" eventid="7788" heatid="25936" lane="2" />
                <ENTRY entrytime="00:00:37.27" eventid="7809" heatid="25952" lane="1" />
                <ENTRY entrytime="00:02:08.60" eventid="1195" heatid="25996" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="26099" firstname="Simone" gender="F" lastname="Aschenbrenner" nation="GER">
              <CONTACT city="SC Schwandorf" />
            </OFFICIAL>
            <OFFICIAL officialid="26049" firstname="Günter" gender="M" lastname="Probst" nation="GER">
              <CONTACT city="SC Schwandorf" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="5147" nation="GER" region="02" clubid="7911" name="Schwimmgemeinschaft Fürth">
          <CONTACT city="Fürth" email="sg.barbara.nestler@gmx.de" name="Nestler Barbara" phone="73 08 28" street="Im Lottersgarten 22" zip="90766" />
          <ATHLETES>
            <ATHLETE birthdate="2007-12-08" firstname="Philipp" gender="M" lastname="Adler" nation="GER" license="407267" athleteid="24263">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.91" entrycourse="SCM" eventid="5702" heatid="25825" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.76" entrycourse="SCM" eventid="5724" heatid="25856" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.20" entrycourse="SCM" eventid="5740" heatid="25903" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.00" eventid="1189" heatid="25983" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-07-10" firstname="Aidan" gender="M" lastname="Amelong" nation="GER" license="370804" athleteid="25593">
              <ENTRIES>
                <ENTRY entrytime="00:03:18.19" entrycourse="SCM" eventid="1177" status="DNS" heatid="25811" lane="4">
                  <MEETINFO city="Lauf" course="SCM" date="2018-01-20" name="Kreismeisterschaften der Jahrgänge 2010 und älter" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.02" entrycourse="SCM" eventid="5702" status="DNS" heatid="25828" lane="2">
                  <MEETINFO city="Lauf" course="SCM" date="2018-01-20" name="Kreismeisterschaften der Jahrgänge 2010 und älter" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.65" entrycourse="SCM" eventid="1141" status="DNS" heatid="25881" lane="4">
                  <MEETINFO city="Lauf" course="SCM" date="2018-01-20" name="Kreismeisterschaften der Jahrgänge 2010 und älter" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.62" entrycourse="SCM" eventid="7773" status="DNS" heatid="25932" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.26" entrycourse="SCM" eventid="1165" status="DNS" heatid="25969" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.94" entrycourse="SCM" eventid="1189" status="DNS" heatid="25989" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-04-01" firstname="Sina" gender="F" lastname="Amelong" nation="GER" license="378026" athleteid="25600">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.89" entrycourse="SCM" eventid="5728" status="DNS" heatid="25871" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.10" entrycourse="SCM" eventid="5744" status="DNS" heatid="25922" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.00" eventid="7788" status="DNS" heatid="25940" lane="1" />
                <ENTRY entrytime="00:00:58.00" eventid="1123" status="DNS" heatid="25962" lane="3" />
                <ENTRY entrytime="00:01:55.68" entrycourse="LCM" eventid="1195" status="DNS" heatid="25998" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-03-11" name="International Swim Meeting Erlangen 2018" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Sinan" gender="M" lastname="Arpert" nation="GER" license="297748" athleteid="24166">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.00" eventid="1177" heatid="25813" lane="1" />
                <ENTRY entrytime="00:00:43.94" eventid="5724" heatid="25863" lane="1" />
                <ENTRY entrytime="00:01:31.60" eventid="1141" heatid="25885" lane="4" />
                <ENTRY entrytime="00:00:43.47" eventid="1117" heatid="25959" lane="3" />
                <ENTRY entrytime="00:01:19.90" eventid="1189" heatid="25991" lane="3" />
                <ENTRY entrytime="00:01:34.34" eventid="7773" heatid="25935" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Ida" gender="F" lastname="Baier" nation="GER" license="347848" athleteid="25304">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.00" eventid="5712" heatid="25845" lane="4" />
                <ENTRY entrytime="00:00:48.07" eventid="5728" heatid="25875" lane="3" />
                <ENTRY entrytime="00:00:40.91" eventid="5744" heatid="25925" lane="5" />
                <ENTRY entrytime="00:01:45.00" eventid="7788" heatid="25943" lane="4" />
                <ENTRY entrytime="00:00:40.00" eventid="1123" heatid="25966" lane="2" />
                <ENTRY entrytime="00:01:37.00" eventid="1195" heatid="26001" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lara" gender="F" lastname="Bamberger" nation="GER" license="362930" athleteid="25455">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.87" eventid="1171" heatid="25976" lane="3" />
                <ENTRY entrytime="00:01:44.63" eventid="1195" heatid="26000" lane="5" />
                <ENTRY entrytime="00:00:52.07" eventid="5712" heatid="25844" lane="1" />
                <ENTRY entrytime="00:00:40.25" eventid="5744" heatid="25925" lane="3" />
                <ENTRY entrytime="00:00:47.88" eventid="5728" heatid="25876" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-09-14" firstname="Sebastian" gender="M" lastname="Behring" nation="GER" license="407268" athleteid="24268">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.71" entrycourse="SCM" eventid="5702" heatid="25829" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.88" entrycourse="SCM" eventid="5724" heatid="25854" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.38" entrycourse="SCM" eventid="5740" heatid="25902" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.00" eventid="1141" heatid="25880" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-10" firstname="Max Eric" gender="M" lastname="Besecke" nation="GER" license="406834" athleteid="25606">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.49" entrycourse="SCM" eventid="1053" heatid="25748" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.63" entrycourse="SCM" eventid="5668" heatid="25759" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.98" entrycourse="SCM" eventid="5678" heatid="25769" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.63" entrycourse="SCM" eventid="7691" heatid="25778" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.63" entrycourse="SCM" eventid="7701" heatid="25807" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-02-17" firstname="Benedek" gender="M" lastname="Boha" nation="GER" license="666666" athleteid="25565">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5702" heatid="25821" lane="3" />
                <ENTRY entrytime="NT" eventid="5724" heatid="25853" lane="2" />
                <ENTRY entrytime="NT" eventid="1141" heatid="25878" lane="2" />
                <ENTRY entrytime="NT" eventid="5740" heatid="25898" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-02" firstname="Dina" gender="F" lastname="Boha" nation="GER" license="391813" athleteid="25612">
              <ENTRIES>
                <ENTRY entrytime="00:01:18.49" entrycourse="LCM" eventid="1195" heatid="26005" lane="5">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-06-30" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
                <ENTRY entrytime="00:03:01.24" entrycourse="LCM" eventid="1183" heatid="25819" lane="5">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-06-30" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.70" entrycourse="SCM" eventid="1111" heatid="25851" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.98" entrycourse="SCM" eventid="1135" heatid="25896" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:27.53" entrycourse="SCM" eventid="1171" heatid="25980" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:03:36.03" entrycourse="SCM" eventid="5661" heatid="26010" lane="2">
                  <MEETINFO city="Nürnberg" course="SCM" date="2018-02-25" name="DMS - Bezirksliga Mittelfranken 2018" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-06-15" firstname="Peter" gender="M" lastname="Boha" nation="GER" athleteid="25570">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25745" lane="5" />
                <ENTRY entrytime="NT" eventid="5668" heatid="25758" lane="6" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25766" lane="3" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25788" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-04-17" firstname="Daniel" gender="M" lastname="Bramigk" nation="GER" license="999999" athleteid="24273">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="5702" heatid="25828" lane="4" />
                <ENTRY entrytime="00:01:02.54" entrycourse="SCM" eventid="5724" heatid="25855" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:48.72" entrycourse="SCM" eventid="5740" heatid="25904" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.00" eventid="7804" heatid="25947" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-06-16" firstname="Anastasia" gender="F" lastname="Chochlow" nation="GER" license="392745" athleteid="25619">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.36" entrycourse="SCM" eventid="5728" heatid="25872" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.00" eventid="5744" heatid="25923" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="7788" heatid="25940" lane="6" />
                <ENTRY entrytime="00:00:48.95" eventid="1123" heatid="25964" lane="4" />
                <ENTRY entrytime="00:01:50.55" eventid="1171" heatid="25977" lane="1" />
                <ENTRY entrytime="00:01:43.41" eventid="1195" heatid="26000" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lena" gender="F" lastname="Clausen" nation="GER" license="99999" athleteid="24208">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5712" heatid="25839" lane="2" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25868" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25917" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Helena" gender="F" lastname="Dautermann" nation="GER" license="393633" athleteid="25311">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.00" eventid="5712" heatid="25846" lane="5" />
                <ENTRY entrytime="00:00:57.11" eventid="5728" heatid="25871" lane="1" />
                <ENTRY entrytime="00:01:50.00" eventid="1135" heatid="25894" lane="3" />
                <ENTRY entrytime="00:00:42.00" eventid="5744" heatid="25924" lane="4" />
                <ENTRY entrytime="00:01:47.00" eventid="1195" heatid="25999" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Simon" gender="M" lastname="Dieret" nation="GER" license="331161" athleteid="24118">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.62" eventid="5724" heatid="25862" lane="3" />
                <ENTRY entrytime="00:00:35.24" eventid="5740" heatid="25911" lane="1" />
                <ENTRY entrytime="00:01:31.68" eventid="7773" heatid="25935" lane="2" />
                <ENTRY entrytime="00:00:41.54" eventid="1117" heatid="25960" lane="1" />
                <ENTRY entrytime="00:01:21.31" eventid="1189" heatid="25991" lane="2" />
                <ENTRY entrytime="00:00:52.92" eventid="5702" heatid="25829" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-04-02" firstname="Leila" gender="F" lastname="Dörrer" nation="GER" license="99999" athleteid="24247">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5664" heatid="25751" lane="4" />
                <ENTRY entrytime="00:01:10.00" eventid="5690" heatid="25795" lane="6" />
                <ENTRY entrytime="00:01:20.00" eventid="7696" heatid="25783" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Alexander" gender="M" lastname="Ehnis" nation="GER" license="331163" athleteid="24173">
              <ENTRIES>
                <ENTRY entrytime="00:02:41.66" eventid="1177" heatid="25813" lane="4" />
                <ENTRY entrytime="00:00:46.73" eventid="5702" heatid="25832" lane="1" />
                <ENTRY entrytime="00:00:33.66" eventid="5740" heatid="25911" lane="4" />
                <ENTRY entrytime="00:01:21.45" eventid="1165" heatid="25972" lane="4" />
                <ENTRY entrytime="00:00:39.44" eventid="5724" heatid="25863" lane="4" />
                <ENTRY entrytime="00:01:13.42" eventid="1189" heatid="25992" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-09-06" firstname="Daniel" gender="M" lastname="Ehnis" nation="GER" license="378024" athleteid="25626">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.00" eventid="1189" heatid="25982" lane="3" />
                <ENTRY entrytime="00:01:04.17" entrycourse="SCM" eventid="5702" heatid="25824" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:08.08" entrycourse="SCM" eventid="5724" heatid="25854" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:05.95" entrycourse="SCM" eventid="5740" heatid="25900" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.00" eventid="7804" heatid="25948" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-09-15" firstname="Julia" gender="F" lastname="Ehnis" nation="GER" athleteid="25632">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.13" entrycourse="SCM" eventid="5664" heatid="25751" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="5674" heatid="25762" lane="3" />
                <ENTRY entrytime="00:01:01.37" entrycourse="SCM" eventid="5682" heatid="25770" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="5690" heatid="25793" lane="3" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25803" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lillian" gender="F" lastname="Ermann" nation="GER" license="279343" athleteid="24125">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.72" eventid="5712" heatid="25847" lane="2" />
                <ENTRY entrytime="00:01:37.81" eventid="1135" heatid="25897" lane="2" />
                <ENTRY entrytime="00:00:40.57" eventid="1123" heatid="25966" lane="5" />
                <ENTRY entrytime="00:01:32.88" eventid="1171" heatid="25979" lane="3" />
                <ENTRY entrytime="00:03:18.60" eventid="5661" heatid="26011" lane="1" />
                <ENTRY entrytime="00:01:28.81" eventid="7788" heatid="25945" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Janis" gender="M" lastname="Fleischmann" nation="GER" license="279338" athleteid="24132">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.28" eventid="1117" heatid="25960" lane="3" />
                <ENTRY entrytime="00:01:13.41" eventid="1165" heatid="25972" lane="3" />
                <ENTRY entrytime="00:01:03.71" eventid="1189" heatid="25992" lane="3" />
                <ENTRY entrytime="00:01:24.53" eventid="1141" heatid="25885" lane="3" />
                <ENTRY entrytime="00:01:12.40" eventid="7773" heatid="25935" lane="3" />
                <ENTRY entrytime="00:00:33.75" eventid="5724" heatid="25863" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-02-15" firstname="Jakob" gender="M" lastname="Freund" nation="GER" license="331165" athleteid="24278">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.69" entrycourse="LCM" eventid="5702" heatid="25827" lane="2">
                  <MEETINFO city="Schwandorf" course="LCM" date="2018-05-12" name="4. Schwandorfer Pokalschwimmfest" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.38" entrycourse="LCM" eventid="1141" heatid="25880" lane="1">
                  <MEETINFO city="Schwandorf" course="LCM" date="2018-05-12" name="4. Schwandorfer Pokalschwimmfest" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.76" entrycourse="SCM" eventid="5740" heatid="25901" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.45" entrycourse="LCM" eventid="1117" heatid="25957" lane="6">
                  <MEETINFO city="Schwandorf" course="LCM" date="2018-05-12" name="4. Schwandorfer Pokalschwimmfest" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-07-11" firstname="Ella Helene" gender="F" lastname="Friedrich" nation="GER" athleteid="25248">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.00" eventid="5674" heatid="25763" lane="2" />
                <ENTRY entrytime="00:00:47.00" eventid="5682" heatid="25771" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" heatid="25784" lane="4" />
                <ENTRY entrytime="00:00:49.00" eventid="5698" heatid="25804" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Anna" gender="F" lastname="Fuchs" nation="GER" license="346281" athleteid="25317">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.00" eventid="5712" heatid="25845" lane="2" />
                <ENTRY entrytime="00:00:49.00" eventid="5728" heatid="25875" lane="5" />
                <ENTRY entrytime="00:00:42.00" eventid="5744" heatid="25924" lane="3" />
                <ENTRY entrytime="00:01:54.00" eventid="7788" heatid="25941" lane="5" />
                <ENTRY entrytime="00:00:24.00" eventid="7809" heatid="25954" lane="2" />
                <ENTRY entrytime="00:01:47.00" eventid="1135" heatid="25895" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lia Sophie" gender="F" lastname="Fuchs" nation="GER" license="0" athleteid="25505">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.65" eventid="5664" heatid="25752" lane="1" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25763" lane="6" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25782" lane="6" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25802" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Maximilian" gender="M" lastname="Fuchs" nation="GER" license="342442" athleteid="25324">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.00" eventid="5702" heatid="25832" lane="6" />
                <ENTRY entrytime="00:01:47.54" eventid="1141" heatid="25884" lane="1" />
                <ENTRY entrytime="00:00:39.79" eventid="5740" heatid="25909" lane="3" />
                <ENTRY entrytime="00:01:55.00" eventid="7773" heatid="25932" lane="4" />
                <ENTRY entrytime="00:01:39.57" eventid="1189" heatid="25988" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Johanna" gender="F" lastname="Geier" nation="GER" license="407274" athleteid="25330">
              <ENTRIES>
                <ENTRY entrytime="00:01:16.46" eventid="5712" heatid="25834" lane="4" />
                <ENTRY entrytime="00:01:15.03" eventid="5728" heatid="25865" lane="3" />
                <ENTRY entrytime="00:01:19.83" eventid="5744" status="DNS" heatid="25914" lane="6" />
                <ENTRY entrytime="00:02:28.00" eventid="1195" heatid="25994" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Roman" gender="M" lastname="Geier" nation="GER" license="347846" athleteid="25335">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.51" eventid="5702" heatid="25831" lane="1" />
                <ENTRY entrytime="00:00:50.77" eventid="5724" heatid="25861" lane="6" />
                <ENTRY entrytime="00:00:48.44" eventid="5740" heatid="25905" lane="6" />
                <ENTRY entrytime="00:01:41.00" eventid="1189" heatid="25987" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="1141" heatid="25883" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jule" gender="F" lastname="Glößinger" nation="GER" license="362932" athleteid="25461">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.09" eventid="5728" heatid="25871" lane="3" />
                <ENTRY entrytime="00:03:56.49" eventid="1183" heatid="25816" lane="2" />
                <ENTRY entrytime="00:01:55.19" eventid="1195" heatid="25998" lane="5" />
                <ENTRY entrytime="00:00:46.20" eventid="5744" heatid="25923" lane="1" />
                <ENTRY entrytime="00:00:56.10" eventid="1123" heatid="25963" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Linnea Emilia" gender="F" lastname="Glößinger" nation="GER" license="389377" athleteid="25510">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.16" eventid="5664" heatid="25753" lane="6" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25782" lane="5" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25793" lane="5" />
                <ENTRY entrytime="00:00:51.91" eventid="5698" heatid="25803" lane="3" />
                <ENTRY entrytime="NT" eventid="7706" heatid="25808" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-06-05" firstname="Philipp" gender="M" lastname="Gorbunov" nation="GER" license="378028" athleteid="25638">
              <ENTRIES>
                <ENTRY entrytime="00:03:59.87" entrycourse="LCM" eventid="1177" heatid="25810" lane="5">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-05-13" name="Erlanger Sparkassen-Cup 2018" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.30" entrycourse="SCM" eventid="5724" heatid="25857" lane="2">
                  <MEETINFO city="Lauf" course="SCM" date="2018-01-20" name="Kreismeisterschaften der Jahrgänge 2010 und älter" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.86" entrycourse="SCM" eventid="5740" heatid="25903" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.00" eventid="1165" heatid="25968" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25985" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-11-12" firstname="Anton" gender="M" lastname="Grießinger" nation="GER" license="362946" athleteid="25644">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.07" entrycourse="LCM" eventid="1177" heatid="25813" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-06-30" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
                <ENTRY entrytime="00:01:39.60" entrycourse="SCM" eventid="1103" heatid="25848" lane="4">
                  <MEETINFO city="Nürnberg" course="SCM" date="2018-02-25" name="DMS - Bezirksliga Mittelfranken 2018" />
                </ENTRY>
                <ENTRY entrytime="00:00:41.26" entrycourse="LCM" eventid="1117" heatid="25960" lane="5">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-07-01" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.62" entrycourse="LCM" eventid="1165" heatid="25972" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-07-01" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
                <ENTRY entrytime="00:01:21.11" entrycourse="SCM" eventid="1189" heatid="25991" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:03:21.53" entrycourse="LCM" eventid="5655" heatid="26007" lane="5">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-07-01" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-02-03" firstname="Peter" gender="M" lastname="Grießinger" nation="GER" license="377882" athleteid="25651">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.23" entrycourse="SCM" eventid="5702" heatid="25827" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:50.91" entrycourse="SCM" eventid="5724" heatid="25860" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.00" eventid="1141" heatid="25883" lane="5" />
                <ENTRY entrytime="NT" eventid="7773" heatid="25929" lane="2" />
                <ENTRY entrytime="NT" eventid="1117" heatid="25956" lane="5" />
                <ENTRY entrytime="00:01:43.00" eventid="1189" heatid="25987" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Levend" gender="M" lastname="Gülec" nation="GER" license="407276" athleteid="25341">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.92" eventid="5702" heatid="25823" lane="3" />
                <ENTRY entrytime="00:01:01.48" eventid="5724" heatid="25855" lane="3" />
                <ENTRY entrytime="00:02:21.00" eventid="1141" heatid="25879" lane="5" />
                <ENTRY entrytime="00:00:54.09" eventid="5740" heatid="25903" lane="1" />
                <ENTRY entrytime="00:02:01.00" eventid="1189" heatid="25983" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Leyan Su" gender="F" lastname="Gülec" nation="GER" license="377883" athleteid="25347">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.66" eventid="5728" heatid="25877" lane="1" />
                <ENTRY entrytime="00:00:36.67" eventid="5744" heatid="25927" lane="3" />
                <ENTRY entrytime="00:01:50.00" eventid="7788" heatid="25942" lane="5" />
                <ENTRY entrytime="00:01:36.47" eventid="1171" heatid="25979" lane="1" />
                <ENTRY entrytime="00:01:32.33" eventid="1195" heatid="26002" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lilith" gender="F" lastname="Heidenreich" nation="GER" license="99999" athleteid="24212">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.00" eventid="5712" heatid="25835" lane="1" />
                <ENTRY entrytime="00:01:30.00" eventid="5744" heatid="25913" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Louisa" gender="F" lastname="Heidenreich" nation="GER" license="99999" athleteid="24215">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.00" eventid="5664" heatid="25752" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="7696" heatid="25783" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="5690" heatid="25795" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Lorena" gender="F" lastname="Heinl" nation="GER" license="407278" athleteid="25353">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.57" eventid="5712" heatid="25842" lane="1" />
                <ENTRY entrytime="00:01:18.75" eventid="5728" heatid="25865" lane="4" />
                <ENTRY entrytime="00:02:40.00" eventid="1135" heatid="25888" lane="4" />
                <ENTRY entrytime="00:00:56.53" eventid="5744" heatid="25918" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-02-21" firstname="Luisa" gender="F" lastname="Heyert" nation="GER" license="347335" athleteid="25658">
              <ENTRIES>
                <ENTRY entrytime="00:03:14.16" entrycourse="SCM" eventid="1183" status="DNS" heatid="25818" lane="2">
                  <MEETINFO city="Nürnberg" course="SCM" date="2018-02-25" name="DMS - Bezirksliga Mittelfranken 2018" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.78" entrycourse="SCM" eventid="1111" status="DNS" heatid="25850" lane="5">
                  <MEETINFO city="Nürnberg" course="SCM" date="2018-02-25" name="DMS - Bezirksliga Mittelfranken 2018" />
                </ENTRY>
                <ENTRY entrytime="00:01:36.68" entrycourse="SCM" eventid="7788" status="DNS" heatid="25944" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:34.02" entrycourse="SCM" eventid="1171" status="DNS" heatid="25979" lane="2">
                  <MEETINFO city="Lauf" course="SCM" date="2018-01-20" name="Kreismeisterschaften der Jahrgänge 2010 und älter" />
                </ENTRY>
                <ENTRY entrytime="00:01:28.99" entrycourse="SCM" eventid="1195" status="DNS" heatid="26003" lane="5">
                  <MEETINFO city="Lauf" course="SCM" date="2018-01-20" name="Kreismeisterschaften der Jahrgänge 2010 und älter" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="5661" status="DNS" heatid="26008" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Tobias" gender="M" lastname="Heyert" nation="GER" license="306630" athleteid="24180">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.11" eventid="5702" heatid="25832" lane="4" />
                <ENTRY entrytime="00:00:33.24" eventid="5740" heatid="25911" lane="3" />
                <ENTRY entrytime="00:00:42.56" eventid="1117" heatid="25960" lane="6" />
                <ENTRY entrytime="00:01:23.53" eventid="1165" heatid="25972" lane="2" />
                <ENTRY entrytime="00:03:08.03" eventid="5655" heatid="26007" lane="3" />
                <ENTRY entrytime="00:02:39.98" eventid="1177" heatid="25813" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Lilly" gender="F" lastname="Hofmann" nation="GER" license="347339" athleteid="24187">
              <ENTRIES>
                <ENTRY entrytime="00:01:24.44" eventid="1111" heatid="25851" lane="3" />
                <ENTRY entrytime="00:00:32.01" eventid="5744" heatid="25928" lane="3" />
                <ENTRY entrytime="00:01:20.65" eventid="1171" heatid="25980" lane="2" />
                <ENTRY entrytime="00:02:53.86" eventid="5661" heatid="26011" lane="3" />
                <ENTRY entrytime="00:02:40.93" eventid="1183" heatid="25820" lane="4" />
                <ENTRY entrytime="00:01:21.53" eventid="7788" heatid="25945" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-08-15" firstname="Sonja" gender="F" lastname="Ilic" nation="GER" license="391815" athleteid="24283">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.91" entrycourse="SCM" eventid="5712" heatid="25839" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:06.43" entrycourse="SCM" eventid="5728" heatid="25867" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.55" entrycourse="SCM" eventid="5744" heatid="25919" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:04.97" entrycourse="SCM" eventid="1123" heatid="25962" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-05" firstname="Emil" gender="M" lastname="Jeske" nation="GER" license="378027" athleteid="25665">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.04" entrycourse="SCM" eventid="5724" heatid="25860" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.61" entrycourse="SCM" eventid="5740" heatid="25909" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="7773" heatid="25930" lane="2" />
                <ENTRY entrytime="NT" eventid="1117" heatid="25956" lane="2" />
                <ENTRY entrytime="00:01:49.13" entrycourse="LCM" eventid="1165" heatid="25970" lane="1">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-03-10" name="International Swim Meeting Erlangen 2018" />
                </ENTRY>
                <ENTRY entrytime="00:01:35.69" entrycourse="LCM" eventid="1189" heatid="25988" lane="2">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-05-13" name="Erlanger Sparkassen-Cup 2018" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Vanessa" gender="F" lastname="Kenner" nation="GER" license="362937" athleteid="25467">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1183" heatid="25814" lane="3" />
                <ENTRY entrytime="00:00:58.95" eventid="5728" heatid="25870" lane="2" />
                <ENTRY entrytime="00:00:49.37" eventid="5744" heatid="25921" lane="5" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25951" lane="2" />
                <ENTRY entrytime="00:02:04.97" eventid="1171" heatid="25975" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Max" gender="M" lastname="Keyser" nation="GER" license="9999" athleteid="24139">
              <ENTRIES>
                <ENTRY entrytime="00:03:30.00" eventid="1177" heatid="25811" lane="6" />
                <ENTRY entrytime="00:00:46.92" eventid="5724" heatid="25862" lane="5" />
                <ENTRY entrytime="00:00:35.63" eventid="5740" heatid="25911" lane="6" />
                <ENTRY entrytime="00:01:35.00" eventid="1189" heatid="25989" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-07-29" firstname="Ferdinand Theo" gender="M" lastname="Krupka" nation="GER" license="99999" athleteid="26012">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" late="yes" heatid="25744" lane="1" />
                <ENTRY entrytime="NT" eventid="7691" late="yes" heatid="25775" lane="4" />
                <ENTRY entrytime="NT" eventid="5686" late="yes" heatid="25786" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-12-16" firstname="Elias" gender="M" lastname="Kunz" nation="GER" license="406835" athleteid="25672">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.81" entrycourse="SCM" eventid="5702" status="DNS" heatid="25823" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.56" entrycourse="SCM" eventid="5724" status="DNS" heatid="25853" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:25.73" entrycourse="SCM" eventid="5740" status="DNS" heatid="25899" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Luca" gender="M" lastname="Lautenschlager" nation="GER" license="404302" athleteid="24308">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.50" eventid="1053" heatid="25747" lane="2" />
                <ENTRY entrytime="00:01:10.00" eventid="5668" heatid="25758" lane="1" />
                <ENTRY entrytime="00:01:10.00" eventid="7691" heatid="25777" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25790" lane="6" />
                <ENTRY entrytime="00:01:05.00" eventid="5694" heatid="25799" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Nils" gender="M" lastname="Lautenschlager" nation="GER" license="372637" athleteid="24314">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.26" eventid="5702" heatid="25823" lane="2" />
                <ENTRY entrytime="00:01:20.82" eventid="5724" heatid="25853" lane="3" />
                <ENTRY entrytime="00:02:30.00" eventid="1141" heatid="25879" lane="1" />
                <ENTRY entrytime="00:01:17.00" eventid="5740" heatid="25900" lane="6" />
                <ENTRY entrytime="00:02:00.00" eventid="1165" status="DNS" heatid="25968" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-06-27" firstname="Edwin" gender="M" lastname="Lichtenwald" nation="GER" license="99999" athleteid="24251">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1053" heatid="25745" lane="3" />
                <ENTRY entrytime="00:01:10.00" eventid="7691" heatid="25777" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25790" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-26" firstname="Livia" gender="F" lastname="Lichtenwald" nation="GER" license="393386" athleteid="25676">
              <ENTRIES>
                <ENTRY entrytime="00:03:48.53" entrycourse="LCM" eventid="1183" heatid="25817" lane="6">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-05-13" name="Erlanger Sparkassen-Cup 2018" />
                </ENTRY>
                <ENTRY entrytime="00:01:58.00" eventid="1135" heatid="25892" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="7788" heatid="25940" lane="5" />
                <ENTRY entrytime="00:00:59.73" entrycourse="SCM" eventid="1123" heatid="25962" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.00" eventid="1195" heatid="26000" lane="6" />
                <ENTRY entrytime="00:01:02.00" eventid="1171" heatid="25980" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Finn" gender="M" lastname="Martin" nation="GER" license="355301" athleteid="25473">
              <ENTRIES>
                <ENTRY entrytime="00:03:11.91" eventid="1177" heatid="25812" lane="1" />
                <ENTRY entrytime="00:01:25.72" eventid="1189" heatid="25990" lane="2" />
                <ENTRY entrytime="00:00:46.29" eventid="5724" heatid="25862" lane="4" />
                <ENTRY entrytime="00:00:36.91" eventid="5740" heatid="25910" lane="2" />
                <ENTRY entrytime="00:01:44.27" eventid="1165" heatid="25970" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Ida" gender="F" lastname="Martin" nation="GER" license="362939" athleteid="25479">
              <ENTRIES>
                <ENTRY entrytime="00:04:11.81" eventid="1183" heatid="25816" lane="6" />
                <ENTRY entrytime="00:01:44.89" eventid="1195" heatid="26000" lane="1" />
                <ENTRY entrytime="00:00:55.66" eventid="5728" heatid="25871" lane="4" />
                <ENTRY entrytime="00:00:48.09" eventid="5744" heatid="25922" lane="6" />
                <ENTRY entrytime="00:00:29.08" eventid="7809" heatid="25952" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Lasse" gender="M" lastname="Martin" nation="GER" license="416998" athleteid="25516">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.59" eventid="1053" status="DNS" heatid="25746" lane="5" />
                <ENTRY entrytime="NT" eventid="5668" status="DNS" heatid="25756" lane="2" />
                <ENTRY entrytime="NT" eventid="7691" status="DNS" heatid="25776" lane="6" />
                <ENTRY entrytime="NT" eventid="5694" status="DNS" heatid="25798" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Nikolaos" gender="M" lastname="Melissourgos" nation="GER" license="365061" athleteid="24144">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.17" eventid="5702" heatid="25830" lane="5" />
                <ENTRY entrytime="00:01:53.53" eventid="1141" heatid="25882" lane="4" />
                <ENTRY entrytime="00:01:45.00" eventid="7773" heatid="25933" lane="3" />
                <ENTRY entrytime="00:00:45.65" eventid="1117" heatid="25959" lane="4" />
                <ENTRY entrytime="00:01:33.92" eventid="1189" heatid="25989" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="David" gender="M" lastname="Milman" nation="GER" license="99999" athleteid="24219">
              <ENTRIES>
                <ENTRY entrytime="00:01:25.00" eventid="5702" heatid="25822" lane="1" />
                <ENTRY entrytime="00:01:30.00" eventid="5740" heatid="25899" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Cosima" gender="F" lastname="Nahr" nation="GER" license="376904" athleteid="24320">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.21" eventid="5712" heatid="25842" lane="3" />
                <ENTRY entrytime="00:01:03.21" eventid="5728" heatid="25869" lane="5" />
                <ENTRY entrytime="00:02:20.00" eventid="1135" heatid="25889" lane="2" />
                <ENTRY entrytime="00:00:55.95" eventid="5744" heatid="25918" lane="4" />
                <ENTRY entrytime="00:02:12.83" eventid="1171" heatid="25974" lane="3" />
                <ENTRY entrytime="00:02:15.95" eventid="1195" heatid="25994" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-09-23" firstname="Julius" gender="M" lastname="Nahr" nation="GER" license="416999" athleteid="24255">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.60" eventid="1053" heatid="25745" lane="2" />
                <ENTRY entrytime="00:01:20.00" eventid="7691" heatid="25776" lane="3" />
                <ENTRY entrytime="00:01:20.00" eventid="5686" heatid="25789" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Maximilian" gender="M" lastname="Neugebauer" nation="GER" license="99999" athleteid="24222">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5724" heatid="25856" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25880" lane="4" />
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25985" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-06-06" firstname="Juliane" gender="F" lastname="Ott" nation="GER" athleteid="25244">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5712" heatid="25837" lane="4" />
                <ENTRY entrytime="00:01:10.00" eventid="5728" heatid="25866" lane="2" />
                <ENTRY entrytime="00:01:05.00" eventid="5744" heatid="25915" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jonas" gender="M" lastname="Penz" nation="GER" license="392570" athleteid="25485">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.53" eventid="5724" heatid="25859" lane="3" />
                <ENTRY entrytime="NT" eventid="1165" heatid="25967" lane="5" />
                <ENTRY entrytime="00:02:02.44" eventid="1189" heatid="25983" lane="2" />
                <ENTRY entrytime="NT" eventid="1177" heatid="25810" lane="6" />
                <ENTRY entrytime="00:00:47.62" eventid="5740" heatid="25905" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Lara" gender="F" lastname="Penz" nation="GER" license="362938" athleteid="25491">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1183" heatid="25814" lane="2" />
                <ENTRY entrytime="00:00:52.27" eventid="5728" heatid="25873" lane="2" />
                <ENTRY entrytime="00:00:39.65" eventid="5744" heatid="25926" lane="6" />
                <ENTRY entrytime="00:00:47.81" eventid="1123" heatid="25965" lane="6" />
                <ENTRY entrytime="NT" eventid="5661" heatid="26008" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-13" firstname="Laurenz" gender="M" lastname="Raum" nation="GER" license="392567" athleteid="25253">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5702" heatid="25824" lane="1" />
                <ENTRY entrytime="00:01:20.00" eventid="5724" heatid="25854" lane="6" />
                <ENTRY entrytime="00:01:05.00" eventid="5740" heatid="25901" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Valentina" gender="F" lastname="Raum" nation="GER" license="337688" athleteid="24150">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.89" eventid="5712" heatid="25846" lane="4" />
                <ENTRY entrytime="00:01:51.65" eventid="1135" heatid="25894" lane="1" />
                <ENTRY entrytime="00:01:43.11" eventid="7788" heatid="25944" lane="1" />
                <ENTRY entrytime="00:00:43.00" eventid="1123" heatid="25966" lane="6" />
                <ENTRY entrytime="00:00:47.85" eventid="5728" heatid="25876" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-12-06" firstname="Clara-Marie" gender="F" lastname="Remiger" nation="GER" license="335471" athleteid="25268">
              <ENTRIES>
                <ENTRY entrytime="00:01:41.33" entrycourse="SCM" eventid="1135" heatid="25896" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2017-06-24" name="16. Bamberg Open 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.66" entrycourse="SCM" eventid="5744" heatid="25926" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.79" entrycourse="SCM" eventid="1123" heatid="25964" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-05-10" firstname="Lian" gender="M" lastname="Richter" nation="GER" license="406841" athleteid="25683">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.95" entrycourse="SCM" eventid="1053" heatid="25749" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.26" entrycourse="SCM" eventid="5668" heatid="25760" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.70" entrycourse="SCM" eventid="5678" heatid="25769" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:38.26" entrycourse="SCM" eventid="7691" heatid="25779" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.14" entrycourse="SCM" eventid="5694" heatid="25801" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-06-22" firstname="Lisa" gender="F" lastname="Rischbeck" nation="GER" license="666666" athleteid="25575">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25750" lane="1" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25763" lane="1" />
                <ENTRY entrytime="NT" eventid="5682" heatid="25770" lane="5" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25783" lane="1" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25803" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-11-12" firstname="THeo" gender="M" lastname="Rischbeck" nation="GER" license="666666" athleteid="25581">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25744" lane="5" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25765" lane="3" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25775" lane="5" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25789" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-06-12" firstname="Sarah-Judith" gender="F" lastname="Ritschke" nation="GER" license="331343" athleteid="25272">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.93" entrycourse="SCM" eventid="5712" heatid="25843" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.72" entrycourse="SCM" eventid="5728" heatid="25873" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.32" entrycourse="SCM" eventid="7788" heatid="25941" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Dennis" gender="M" lastname="Rosenthal" nation="GER" license="347337" athleteid="24156">
              <ENTRIES>
                <ENTRY entrytime="00:03:24.22" eventid="1177" heatid="25811" lane="1" />
                <ENTRY entrytime="00:00:49.01" eventid="5724" heatid="25861" lane="4" />
                <ENTRY entrytime="00:00:39.56" eventid="5740" heatid="25910" lane="6" />
                <ENTRY entrytime="00:01:33.47" eventid="1189" heatid="25989" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Frank" gender="M" lastname="Rosenthal" nation="GER" athleteid="24327">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="1053" heatid="25746" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5668" heatid="25758" lane="2" />
                <ENTRY entrytime="00:01:00.00" eventid="5686" heatid="25790" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Robin" gender="M" lastname="Rosenthal" nation="GER" license="362942" athleteid="25358">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.80" eventid="5702" heatid="25827" lane="1" />
                <ENTRY entrytime="00:02:16.52" eventid="1141" heatid="25879" lane="3" />
                <ENTRY entrytime="00:01:07.56" eventid="1117" heatid="25956" lane="4" />
                <ENTRY entrytime="00:01:57.77" eventid="1189" heatid="25984" lane="2" />
                <ENTRY entrytime="00:02:09.00" eventid="7773" heatid="25931" lane="5" />
                <ENTRY entrytime="00:01:57.00" eventid="1165" heatid="25969" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-07-10" firstname="Ronja" gender="F" lastname="Rosenthal" nation="GER" license="389376" athleteid="25689">
              <ENTRIES>
                <ENTRY entrytime="00:03:45.00" eventid="1183" heatid="25817" lane="1" />
                <ENTRY entrytime="00:00:56.65" entrycourse="SCM" eventid="5728" heatid="25871" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:59.00" eventid="1135" heatid="25892" lane="5" />
                <ENTRY entrytime="00:00:49.00" eventid="5744" heatid="25921" lane="3" />
                <ENTRY entrytime="00:02:00.00" eventid="1171" heatid="25976" lane="1" />
                <ENTRY entrytime="00:01:58.00" eventid="1195" heatid="25997" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Leana Isabel" gender="F" lastname="Rother" nation="GER" license="379366" athleteid="24331">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.54" eventid="5712" heatid="25842" lane="5" />
                <ENTRY entrytime="00:01:01.24" eventid="5728" heatid="25870" lane="6" />
                <ENTRY entrytime="00:02:20.00" eventid="1135" heatid="25889" lane="4" />
                <ENTRY entrytime="00:00:51.03" eventid="5744" heatid="25920" lane="2" />
                <ENTRY entrytime="00:02:30.00" eventid="1195" heatid="25993" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Timon Sebastian" gender="M" lastname="Rother" nation="GER" license="406840" athleteid="24337">
              <ENTRIES>
                <ENTRY entrytime="00:00:38.70" eventid="1053" heatid="25747" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5668" heatid="25758" lane="5" />
                <ENTRY entrytime="00:01:10.00" eventid="7691" heatid="25777" lane="5" />
                <ENTRY entrytime="00:01:10.00" eventid="5686" heatid="25789" lane="3" />
                <ENTRY entrytime="00:00:44.61" eventid="5678" heatid="25767" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Erem Sonsuz" gender="M" lastname="Sahin" nation="GER" license="378025" athleteid="25365">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.98" eventid="5702" heatid="25830" lane="2" />
                <ENTRY entrytime="00:00:59.00" eventid="5724" heatid="25856" lane="3" />
                <ENTRY entrytime="00:01:53.58" eventid="1141" heatid="25882" lane="5" />
                <ENTRY entrytime="00:00:49.00" eventid="5740" heatid="25904" lane="5" />
                <ENTRY entrytime="00:01:43.00" eventid="1189" heatid="25986" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-05-03" firstname="Elina" gender="F" lastname="Sandig" nation="GER" license="392573" athleteid="25257">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.54" entrycourse="SCM" eventid="5664" heatid="25754" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.00" eventid="5674" heatid="25763" lane="3" />
                <ENTRY entrytime="00:00:31.92" entrycourse="SCM" eventid="5682" heatid="25773" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.00" eventid="5690" heatid="25796" lane="2" />
                <ENTRY entrytime="00:00:35.06" entrycourse="SCM" eventid="5698" heatid="25805" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Jonathan" gender="M" lastname="Sandig" nation="GER" license="413757" athleteid="25497">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5702" heatid="25822" lane="6" />
                <ENTRY entrytime="NT" eventid="5724" heatid="25852" lane="2" />
                <ENTRY entrytime="NT" eventid="5740" heatid="25898" lane="2" />
                <ENTRY entrytime="NT" eventid="1189" heatid="25981" lane="2" />
                <ENTRY entrytime="NT" eventid="1165" heatid="25967" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-06-24" firstname="Diana" gender="F" lastname="Satsevich" nation="GER" license="666666" athleteid="25586">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.00" eventid="7788" heatid="25943" lane="2" />
                <ENTRY entrytime="00:01:40.50" eventid="1171" heatid="25978" lane="4" />
                <ENTRY entrytime="00:01:22.50" eventid="1195" heatid="26004" lane="4" />
                <ENTRY entrytime="00:03:02.90" eventid="1183" heatid="25819" lane="1" />
                <ENTRY entrytime="00:00:52.00" eventid="5712" heatid="25844" lane="5" />
                <ENTRY entrytime="00:01:52.00" eventid="1135" heatid="25894" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Jan" gender="M" lastname="Schafner" nation="GER" license="406833" athleteid="25521">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.06" eventid="1053" heatid="25747" lane="5" />
                <ENTRY entrytime="NT" eventid="5668" heatid="25756" lane="5" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25766" lane="4" />
                <ENTRY entrytime="NT" eventid="7691" heatid="25776" lane="1" />
                <ENTRY entrytime="00:00:42.37" eventid="5694" heatid="25799" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Julian" gender="M" lastname="Schafner" nation="GER" license="359179" athleteid="25371">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.28" eventid="5702" heatid="25831" lane="4" />
                <ENTRY entrytime="00:00:51.31" eventid="5724" heatid="25860" lane="2" />
                <ENTRY entrytime="00:01:42.00" eventid="1141" heatid="25884" lane="4" />
                <ENTRY entrytime="00:00:39.00" eventid="5740" heatid="25910" lane="1" />
                <ENTRY entrytime="00:01:44.00" eventid="7773" heatid="25934" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="1117" heatid="25958" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Clara" gender="F" lastname="Schiller" nation="GER" license="99999" athleteid="24226">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5712" heatid="25837" lane="3" />
                <ENTRY entrytime="00:01:05.00" eventid="5744" heatid="25915" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Elsa" gender="F" lastname="Schmaus" nation="GER" license="99999" athleteid="24229">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="5698" heatid="25803" lane="4" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" heatid="25784" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Greta" gender="F" lastname="Schmaus" nation="GER" license="403439" athleteid="25378">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.84" eventid="5712" heatid="25840" lane="3" />
                <ENTRY entrytime="00:00:58.94" eventid="5728" heatid="25870" lane="4" />
                <ENTRY entrytime="00:02:10.58" eventid="1135" heatid="25890" lane="3" />
                <ENTRY entrytime="00:00:54.48" eventid="5744" heatid="25919" lane="2" />
                <ENTRY entrytime="00:01:58.00" eventid="1195" heatid="25997" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Finja" gender="F" lastname="Schmidt" nation="GER" license="362945" athleteid="25384">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.00" eventid="5712" heatid="25843" lane="3" />
                <ENTRY entrytime="00:00:48.00" eventid="5728" heatid="25876" lane="6" />
                <ENTRY entrytime="00:00:39.00" eventid="5744" heatid="25926" lane="1" />
                <ENTRY entrytime="00:01:51.00" eventid="7788" heatid="25941" lane="4" />
                <ENTRY entrytime="00:00:23.90" eventid="7809" heatid="25954" lane="3" />
                <ENTRY entrytime="00:01:46.00" eventid="1195" heatid="25999" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Leoni" gender="F" lastname="Schmidt" nation="GER" license="331171" athleteid="25391">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.00" eventid="5712" heatid="25845" lane="6" />
                <ENTRY entrytime="00:00:49.00" eventid="5728" heatid="25875" lane="2" />
                <ENTRY entrytime="00:00:39.00" eventid="5744" heatid="25926" lane="5" />
                <ENTRY entrytime="00:01:50.00" eventid="7788" heatid="25942" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="1123" heatid="25964" lane="6" />
                <ENTRY entrytime="00:01:35.00" eventid="1195" heatid="26002" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-10-27" firstname="Celia Zoé" gender="F" lastname="Schnake" nation="GER" license="385213" athleteid="25696">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.37" entrycourse="SCM" eventid="5712" heatid="25842" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.95" entrycourse="SCM" eventid="5728" heatid="25875" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="25892" lane="6" />
                <ENTRY entrytime="00:00:46.61" entrycourse="SCM" eventid="5744" heatid="25922" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.00" eventid="1195" heatid="25999" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-10-28" firstname="Emily" gender="F" lastname="Schramm" nation="GER" athleteid="25263">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.00" eventid="5674" heatid="25763" lane="4" />
                <ENTRY entrytime="00:00:45.00" eventid="5682" heatid="25771" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" heatid="25784" lane="5" />
                <ENTRY entrytime="00:00:47.00" eventid="5698" heatid="25804" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-02-16" firstname="Lara" gender="F" lastname="Schuler" nation="GER" license="348128" athleteid="25276">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.92" entrycourse="SCM" eventid="5728" heatid="25875" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:47.70" entrycourse="SCM" eventid="1135" heatid="25895" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2017-06-24" name="16. Bamberg Open 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.72" entrycourse="SCM" eventid="5744" heatid="25925" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-11-24" firstname="Luca" gender="M" lastname="Schuler" nation="GER" license="393384" athleteid="25280">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25880" lane="2" />
                <ENTRY entrytime="00:00:47.86" entrycourse="SCM" eventid="5740" heatid="25905" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.00" eventid="7804" heatid="25947" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Cem Leon" gender="M" lastname="Schulze Döring" nation="GER" license="346286" athleteid="24201">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.71" eventid="5702" heatid="25832" lane="2" />
                <ENTRY entrytime="00:00:44.33" eventid="5724" heatid="25863" lane="6" />
                <ENTRY entrytime="00:00:46.41" eventid="1117" heatid="25959" lane="2" />
                <ENTRY entrytime="00:01:18.46" eventid="1189" heatid="25992" lane="6" />
                <ENTRY entrytime="00:03:18.57" eventid="5655" heatid="26007" lane="2" />
                <ENTRY entrytime="00:01:33.43" eventid="7773" heatid="25935" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-24" firstname="Finn Tolgar" gender="M" lastname="Schulze Döring" nation="GER" license="368690" athleteid="25702">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.59" entrycourse="SCM" eventid="1053" heatid="25749" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.92" entrycourse="SCM" eventid="5668" heatid="25760" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.10" entrycourse="SCM" eventid="5678" heatid="25769" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.92" entrycourse="SCM" eventid="7691" heatid="25779" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.68" entrycourse="SCM" eventid="5694" heatid="25801" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-07-30" firstname="Nils Ömer" gender="M" lastname="Schulze Döring" nation="GER" license="393382" athleteid="25708">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.94" entrycourse="SCM" eventid="1053" heatid="25749" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.41" entrycourse="SCM" eventid="5668" heatid="25759" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.15" entrycourse="SCM" eventid="5678" heatid="25769" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.41" entrycourse="SCM" eventid="7691" heatid="25777" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.54" entrycourse="SCM" eventid="5694" heatid="25800" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Antonia" gender="F" lastname="Schödl" nation="GER" athleteid="25527">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25751" lane="6" />
                <ENTRY entrytime="NT" eventid="5674" heatid="25763" lane="5" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25803" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Franziska" gender="F" lastname="Schöttl" nation="GER" license="322657" athleteid="24194">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.48" eventid="5712" heatid="25845" lane="1" />
                <ENTRY entrytime="00:02:00.41" eventid="1111" heatid="25849" lane="2" />
                <ENTRY entrytime="00:00:40.26" eventid="5744" heatid="25925" lane="4" />
                <ENTRY entrytime="00:01:42.34" eventid="1171" heatid="25977" lane="3" />
                <ENTRY entrytime="00:03:51.68" eventid="5661" heatid="26009" lane="5" />
                <ENTRY entrytime="00:01:46.50" eventid="7788" heatid="25943" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-10-01" firstname="Stefan" gender="M" lastname="Schütz" nation="GER" license="368692" athleteid="25284">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.66" entrycourse="SCM" eventid="5702" status="DNS" heatid="25825" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.36" entrycourse="SCM" eventid="1117" status="DNS" heatid="25958" lane="6">
                  <MEETINFO city="Wackersdorf" course="SCM" date="2017-07-15" name="5. Wackersdorfer Panoramabad-Schwimmfest 2017" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.48" entrycourse="SCM" eventid="1189" status="DNS" heatid="25987" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-05-28" firstname="Tamara" gender="F" lastname="Sladojevic" nation="GER" license="378023" athleteid="24288">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.36" entrycourse="SCM" eventid="5712" heatid="25843" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:02.61" entrycourse="SCM" eventid="5728" heatid="25869" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.34" entrycourse="SCM" eventid="5744" heatid="25920" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.00" eventid="1135" heatid="25891" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-03-26" firstname="Tijana" gender="F" lastname="Sladojevic" nation="GER" license="362941" athleteid="24293">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.91" entrycourse="SCM" eventid="5728" heatid="25872" lane="5">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.00" entrycourse="SCM" eventid="5744" heatid="25924" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.00" eventid="1135" heatid="25894" lane="5" />
                <ENTRY entrytime="00:01:55.00" eventid="1171" heatid="25976" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Dominik" gender="M" lastname="Slonicz" nation="GER" license="000000" athleteid="24343">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25744" lane="4" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25786" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2013-01-01" firstname="Julia" gender="F" lastname="Slonicz" nation="GER" license="000000" athleteid="24346">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25751" lane="2" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25792" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-08-10" firstname="Elena" gender="F" lastname="Stoll" nation="GER" license="295232" athleteid="25288">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.30" entrycourse="SCM" eventid="5728" heatid="25876" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.11" entrycourse="SCM" eventid="5744" heatid="25927" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.97" entrycourse="SCM" eventid="7788" heatid="25944" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-08-10" firstname="Nicola" gender="F" lastname="Stoll" nation="GER" license="295233" athleteid="25292">
              <ENTRIES>
                <ENTRY entrytime="00:02:58.27" entrycourse="SCM" eventid="1183" heatid="25819" lane="3">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:36.96" entrycourse="SCM" eventid="5744" heatid="25927" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:44.66" entrycourse="SCM" eventid="1123" heatid="25965" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-25" firstname="Roman" gender="M" lastname="Stroh" nation="GER" license="413758" athleteid="25714">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5702" status="DNS" heatid="25821" lane="1" />
                <ENTRY entrytime="NT" eventid="5724" status="DNS" heatid="25852" lane="4" />
                <ENTRY entrytime="NT" eventid="5740" status="DNS" heatid="25899" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Amir" gender="M" lastname="Tawfik" nation="GER" license="99999" athleteid="24232">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.00" eventid="1053" heatid="25746" lane="1" />
                <ENTRY entrytime="00:00:50.00" eventid="5686" heatid="25790" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Amira" gender="F" lastname="Tawfik" nation="GER" license="99999" athleteid="24235">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.00" eventid="5698" heatid="25804" lane="2" />
                <ENTRY entrytime="00:00:40.00" eventid="5664" heatid="25753" lane="5" />
                <ENTRY entrytime="00:00:50.00" eventid="7696" heatid="25784" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Annika" gender="F" lastname="Thummerer" nation="GER" license="393378" athleteid="25398">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.00" eventid="5712" heatid="25838" lane="2" />
                <ENTRY entrytime="00:01:04.75" eventid="5728" heatid="25868" lane="4" />
                <ENTRY entrytime="00:02:13.00" eventid="1135" heatid="25890" lane="4" />
                <ENTRY entrytime="00:00:59.00" eventid="5744" heatid="25917" lane="4" />
                <ENTRY entrytime="00:02:10.00" eventid="7788" heatid="25939" lane="1" />
                <ENTRY entrytime="00:00:31.00" eventid="7809" heatid="25952" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Carla" gender="F" lastname="Timpe" nation="GER" license="377884" athleteid="25405">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.60" eventid="5712" heatid="25841" lane="6" />
                <ENTRY entrytime="00:01:06.47" eventid="5728" heatid="25867" lane="6" />
                <ENTRY entrytime="00:02:10.33" eventid="1135" heatid="25891" lane="6" />
                <ENTRY entrytime="00:00:49.77" eventid="5744" heatid="25921" lane="6" />
                <ENTRY entrytime="00:01:49.00" eventid="1195" heatid="25999" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Winnie" gender="F" lastname="Waßmuth" nation="GER" athleteid="25531">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25751" lane="5" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25782" lane="2" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25793" lane="4" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25803" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-04" firstname="Emily" gender="F" lastname="Wech" nation="GER" license="359178" athleteid="24298">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.98" entrycourse="SCM" eventid="7788" heatid="25939" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.12" entrycourse="SCM" eventid="1135" heatid="25891" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.92" entrycourse="SCM" eventid="1123" heatid="25963" lane="1">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.96" entrycourse="SCM" eventid="1171" heatid="25975" lane="4">
                  <MEETINFO course="SCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leander" gender="M" lastname="Wech" nation="GER" license="392571" athleteid="24239">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5702" heatid="25823" lane="1" />
                <ENTRY entrytime="00:01:05.00" eventid="5724" heatid="25854" lane="3" />
                <ENTRY entrytime="00:01:05.00" eventid="5740" heatid="25901" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-10-19" firstname="Patrick" gender="M" lastname="Wech" nation="GER" license="392572" athleteid="24303">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.59" entrycourse="SCM" eventid="5702" heatid="25824" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.33" entrycourse="SCM" eventid="5724" heatid="25857" lane="3">
                  <MEETINFO city="Fürth" course="SCM" date="2017-11-11" name="41. Fürther Kinderschwimmen" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.60" entrycourse="SCM" eventid="5740" heatid="25907" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.00" eventid="1165" heatid="25969" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Anna-Lena" gender="F" lastname="Weisbrodt" nation="GER" license="407277" athleteid="25411">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.00" eventid="5712" heatid="25840" lane="6" />
                <ENTRY entrytime="00:01:05.41" eventid="5728" heatid="25867" lane="5" />
                <ENTRY entrytime="00:02:19.00" eventid="1135" heatid="25889" lane="3" />
                <ENTRY entrytime="00:00:53.51" eventid="5744" heatid="25919" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-05-01" firstname="Michael" gender="M" lastname="Wiegandt" nation="GER" license="392893" athleteid="25718">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.89" entrycourse="SCM" eventid="5702" heatid="25830" lane="4">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.20" entrycourse="SCM" eventid="5724" heatid="25859" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:45.31" entrycourse="SCM" eventid="5740" heatid="25907" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="7773" heatid="25929" lane="4" />
                <ENTRY entrytime="00:01:46.83" entrycourse="LCM" eventid="1189" heatid="25986" lane="5">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-05-13" name="Erlanger Sparkassen-Cup 2018" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-05-12" firstname="Lukas" gender="M" lastname="Wildner" nation="GER" license="348129" athleteid="25300">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.00" entrycourse="SCM" eventid="5740" heatid="25908" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.33" entrycourse="SCM" eventid="1117" heatid="25959" lane="6">
                  <MEETINFO city="Fürth" course="SCM" date="2017-03-25" name="SG Fürth Vereinsmeisterschaften 2017" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:23.04" entrycourse="SCM" eventid="1189" heatid="25991" lane="6">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-06-07" firstname="Caspar-Julius" gender="M" lastname="Wilke" nation="GER" license="368701" athleteid="25724">
              <ENTRIES>
                <ENTRY entrytime="00:02:50.98" entrycourse="LCM" eventid="1177" heatid="25813" lane="2">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-06-30" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.44" entrycourse="SCM" eventid="1103" heatid="25848" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.56" entrycourse="SCM" eventid="1141" heatid="25885" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:37.72" entrycourse="SCM" eventid="1165" heatid="25971" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:30.25" eventid="1189" heatid="25981" lane="4" />
                <ENTRY entrytime="00:03:11.46" entrycourse="LCM" eventid="5655" heatid="26007" lane="4">
                  <MEETINFO city="Erlangen" course="LCM" date="2018-07-01" name="Bezirks Jahrgangs- und Juniorenmeisterschaften Mittelfraenkische Meisterschaften" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-01-01" firstname="Annika" gender="F" lastname="Wolf" nation="GER" license="407273" athleteid="24161">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.27" eventid="5712" status="DNS" heatid="25846" lane="2" />
                <ENTRY entrytime="00:00:43.30" eventid="5728" status="DNS" heatid="25877" lane="2" />
                <ENTRY entrytime="00:00:37.54" eventid="5744" status="DNS" heatid="25926" lane="3" />
                <ENTRY entrytime="00:01:30.00" eventid="1195" status="DNS" heatid="26003" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-11-19" firstname="Julia" gender="F" lastname="Wolf" nation="GER" license="362947" athleteid="25731">
              <ENTRIES>
                <ENTRY entrytime="00:03:23.68" entrycourse="SCM" eventid="1183" heatid="25818" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:01:38.13" entrycourse="SCM" eventid="1111" heatid="25850" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.73" entrycourse="SCM" eventid="1135" heatid="25895" lane="3">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.52" entrycourse="SCM" eventid="1171" heatid="25978" lane="5">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:01:29.06" entrycourse="SCM" eventid="1195" heatid="26003" lane="1">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.00" eventid="5661" heatid="26010" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-12-26" firstname="Jan" gender="M" lastname="Zeidler" nation="GER" license="389378" athleteid="25738">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.00" eventid="5686" status="DNS" heatid="25791" lane="2" />
                <ENTRY entrytime="00:00:31.03" entrycourse="SCM" eventid="1053" status="DNS" heatid="25749" lane="6">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.00" eventid="5668" status="DNS" heatid="25760" lane="2" />
                <ENTRY entrytime="00:00:36.99" entrycourse="SCM" eventid="5678" status="DNS" heatid="25768" lane="2">
                  <MEETINFO course="SCM" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.00" eventid="5694" status="DNS" heatid="25800" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2004-09-18" firstname="Tim" gender="M" lastname="Überla" nation="GER" license="331340" athleteid="25296">
              <ENTRIES>
                <ENTRY entrytime="00:01:32.65" entrycourse="SCM" eventid="1141" heatid="25885" lane="2">
                  <MEETINFO city="Bamberg" course="SCM" date="2018-06-16" name="17. Bamberg Open 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.75" entrycourse="SCM" eventid="5740" heatid="25910" lane="4">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.94" entrycourse="SCM" eventid="1117" heatid="25958" lane="2">
                  <MEETINFO city="Fürth" course="SCM" date="2018-01-27" name="SG Fürth Vereinsmeisterschaften 2018" nation="GER" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="8" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="23774" heatid="25946" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="24293" number="1" />
                    <RELAYPOSITION athleteid="25324" number="2" />
                    <RELAYPOSITION athleteid="24298" number="3" />
                    <RELAYPOSITION athleteid="25371" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="26026" firstname="Samuel" gender="M" lastname="Arpert" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26041" firstname="Ulrich" gender="M" lastname="Arpert" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26030" firstname="Henri" gender="M" lastname="Babinsky" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26097" firstname="Daniela" gender="F" lastname="Erdmann" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26096" firstname="Wolfgang" gender="M" lastname="Ermann" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26024" firstname="Matthias" gender="M" lastname="Fuchs" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26045" firstname="Natascha" gender="F" lastname="Griesinger" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26032" firstname="Ruth" gender="F" lastname="Papuschek" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26117" firstname="Roman" gender="M" lastname="Penz" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26039" firstname="Daniel" gender="M" lastname="Pfob" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26037" firstname="Dominikus" gender="M" lastname="Schmitt" nation="GER">
              <CONTACT city="SG Fürth" />
            </OFFICIAL>
            <OFFICIAL officialid="26100" firstname="Richard" gender="M" lastname="Schöttl" nation="GER">
              <CONTACT city="SG Füth" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="5498" nation="GER" region="02" clubid="7947" name="Schwimmgemeinschaft-Lauf">
          <OFFICIALS>
            <OFFICIAL officialid="17218" firstname="Isabel" gender="F" lastname="Goltz" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4301" nation="GER" region="02" clubid="7917" name="Schwimmteam Neusäß" />
        <CLUB type="CLUB" code="4344" nation="GER" region="02" clubid="7930" name="SCHWIMMVEREIN AUGSBURG 1911 e.V." shortname="SCHWIMMVEREIN AUGSBURG 1911 e." />
        <CLUB type="CLUB" code="6399" nation="GER" region="02" clubid="7961" name="SG - Elsenfeld/Kleinwallstadt" />
        <CLUB type="CLUB" code="5085" nation="GER" region="02" clubid="7923" name="SG Bamberg" />
        <CLUB type="CLUB" code="5438" nation="GER" region="02" clubid="7973" name="SG Ergolding/Landau" />
        <CLUB type="CLUB" code="5095" nation="GER" region="02" clubid="7886" name="SG Frankenhöhe">
          <OFFICIALS>
            <OFFICIAL officialid="17201" firstname="Daniela" gender="F" lastname="Gräf" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="5068" nation="GER" region="02" clubid="7896" name="SG Haßberge" />
        <CLUB type="CLUB" code="5212" nation="GER" region="2" clubid="7966" name="SG Mallersdorf/Pfaffenberg" />
        <CLUB type="CLUB" code="6768" nation="GER" region="02" clubid="7945" name="SG Mittelfranken">
          <ATHLETES>
            <ATHLETE birthdate="2006-01-01" firstname="Marco" gender="M" lastname="Arnis" nation="GER" license="371878" athleteid="24708">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.96" eventid="1141" heatid="25884" lane="5" />
                <ENTRY entrytime="00:01:39.80" eventid="7773" heatid="25934" lane="2" />
                <ENTRY entrytime="00:00:50.69" eventid="1117" heatid="25958" lane="4" />
                <ENTRY entrytime="00:01:38.44" eventid="1165" heatid="25971" lane="1" />
                <ENTRY entrytime="00:01:28.37" eventid="1189" heatid="25990" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Paulina" gender="F" lastname="Artavia" nation="GER" license="377714" athleteid="24714">
              <ENTRIES>
                <ENTRY entrytime="00:01:44.25" eventid="1135" heatid="25896" lane="1" />
                <ENTRY entrytime="00:01:34.92" eventid="7788" heatid="25945" lane="5" />
                <ENTRY entrytime="00:00:42.03" eventid="1123" heatid="25966" lane="1" />
                <ENTRY entrytime="00:01:31.60" eventid="1171" heatid="25980" lane="6" />
                <ENTRY entrytime="00:01:30.66" eventid="1195" heatid="26002" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Liv" gender="F" lastname="Asse" nation="GER" license="406748" athleteid="24720">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.56" eventid="5712" heatid="25839" lane="6" />
                <ENTRY entrytime="00:00:53.20" eventid="5728" heatid="25873" lane="5" />
                <ENTRY entrytime="00:00:49.31" eventid="5744" heatid="25921" lane="2" />
                <ENTRY entrytime="00:01:55.00" eventid="7788" heatid="25940" lane="4" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25954" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Martin" gender="M" lastname="Bachmann" nation="GER" license="382799" athleteid="24726">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.04" eventid="5702" heatid="25828" lane="1" />
                <ENTRY entrytime="00:00:54.20" eventid="5724" heatid="25859" lane="1" />
                <ENTRY entrytime="00:00:47.95" eventid="5740" heatid="25905" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Any" gender="F" lastname="Bauer-Makichyan" nation="GER" license="420703" athleteid="25536">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25834" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Anthony" gender="M" lastname="Blumenthal" nation="GER" license="403952" athleteid="25105">
              <ENTRIES>
                <ENTRY entrytime="00:00:41.16" eventid="5724" heatid="25863" lane="2" />
                <ENTRY entrytime="00:00:34.02" eventid="5740" heatid="25911" lane="5" />
                <ENTRY entrytime="00:01:37.31" eventid="7773" heatid="25934" lane="3" />
                <ENTRY entrytime="00:01:26.24" eventid="1165" heatid="25972" lane="1" />
                <ENTRY entrytime="00:01:18.43" eventid="1189" heatid="25992" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Laura" gender="F" lastname="Blumenthal" nation="GER" license="403951" athleteid="25099">
              <ENTRIES>
                <ENTRY entrytime="00:02:54.07" eventid="1183" heatid="25820" lane="6" />
                <ENTRY entrytime="00:00:43.25" eventid="5728" heatid="25877" lane="4" />
                <ENTRY entrytime="00:00:35.23" eventid="5744" heatid="25928" lane="2" />
                <ENTRY entrytime="00:01:32.95" eventid="1171" heatid="25979" lane="4" />
                <ENTRY entrytime="00:01:18.68" eventid="1195" heatid="26005" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Sebastian" gender="M" lastname="Brandner" nation="GER" license="406001" athleteid="24734">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.96" eventid="5702" heatid="25827" lane="6" />
                <ENTRY entrytime="00:00:50.42" eventid="5724" heatid="25861" lane="1" />
                <ENTRY entrytime="00:00:42.00" eventid="5740" heatid="25908" lane="5" />
                <ENTRY entrytime="00:02:05.00" eventid="7773" heatid="25931" lane="4" />
                <ENTRY entrytime="00:00:23.07" eventid="7804" heatid="25949" lane="4" />
                <ENTRY entrytime="00:01:47.92" eventid="1189" heatid="25986" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Pia" gender="F" lastname="Braun" nation="GER" license="383927" athleteid="24741">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.44" eventid="5712" heatid="25846" lane="3" />
                <ENTRY entrytime="00:00:54.00" eventid="5728" heatid="25872" lane="3" />
                <ENTRY entrytime="00:00:42.69" eventid="5744" heatid="25924" lane="2" />
                <ENTRY entrytime="00:02:05.00" eventid="7788" heatid="25939" lane="4" />
                <ENTRY entrytime="00:00:23.00" eventid="7809" heatid="25955" lane="6" />
                <ENTRY entrytime="00:01:44.23" eventid="1195" heatid="26000" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Isabelle Zoe" gender="F" lastname="Brauns" nation="GER" license="415616" athleteid="24748">
              <ENTRIES>
                <ENTRY entrytime="00:02:16.92" eventid="1135" heatid="25890" lane="2" />
                <ENTRY entrytime="00:01:04.19" eventid="5744" heatid="25916" lane="6" />
                <ENTRY entrytime="00:02:10.23" eventid="7788" heatid="25939" lane="6" />
                <ENTRY entrytime="00:02:09.28" eventid="1171" heatid="25975" lane="5" />
                <ENTRY entrytime="00:02:09.32" eventid="1195" heatid="25995" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Leonie Emma" gender="F" lastname="Brauns" nation="GER" license="406688" athleteid="24754">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.73" eventid="5712" heatid="25842" lane="6" />
                <ENTRY entrytime="00:00:51.28" eventid="5728" heatid="25874" lane="1" />
                <ENTRY entrytime="00:02:01.73" eventid="1135" heatid="25891" lane="2" />
                <ENTRY entrytime="00:00:44.85" eventid="5744" heatid="25923" lane="3" />
                <ENTRY entrytime="00:01:47.89" eventid="1171" heatid="25977" lane="5" />
                <ENTRY entrytime="00:01:43.11" eventid="1195" heatid="26000" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Helena" gender="F" lastname="Brausum" nation="GER" license="420240" athleteid="24761">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25836" lane="6" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25867" lane="3" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25917" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Luisa" gender="F" lastname="Brückner" nation="GER" license="416118" athleteid="24765">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.01" eventid="5712" heatid="25838" lane="4" />
                <ENTRY entrytime="00:00:54.82" eventid="5728" heatid="25872" lane="2" />
                <ENTRY entrytime="00:00:46.60" eventid="5744" heatid="25922" lane="3" />
                <ENTRY entrytime="00:01:55.00" eventid="7788" heatid="25941" lane="6" />
                <ENTRY entrytime="00:00:25.75" eventid="7809" heatid="25953" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Paul Wilfried Jens" gender="M" lastname="Burkhardt" nation="GER" license="406751" athleteid="24771">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.46" eventid="5702" heatid="25823" lane="5" />
                <ENTRY entrytime="00:00:55.31" eventid="5724" heatid="25858" lane="5" />
                <ENTRY entrytime="00:00:52.63" eventid="5740" heatid="25903" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Michael" gender="M" lastname="Burla" nation="GER" license="417322" athleteid="24775">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.00" eventid="5702" heatid="25825" lane="4" />
                <ENTRY entrytime="00:00:58.00" eventid="5724" heatid="25857" lane="5" />
                <ENTRY entrytime="00:00:53.00" eventid="5740" heatid="25903" lane="5" />
                <ENTRY entrytime="00:02:15.00" eventid="7773" heatid="25931" lane="6" />
                <ENTRY entrytime="00:00:29.00" eventid="7804" status="DNS" heatid="25948" lane="1" />
                <ENTRY entrytime="00:02:09.00" eventid="1189" heatid="25983" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Chiara" gender="F" lastname="Böller" nation="GER" license="392887" athleteid="24730">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.97" eventid="5728" heatid="25873" lane="3" />
                <ENTRY entrytime="00:01:47.47" eventid="1135" heatid="25895" lane="1" />
                <ENTRY entrytime="00:00:46.36" eventid="5744" heatid="25923" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Sophie" gender="F" lastname="Böller" nation="GER" athleteid="25084">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25836" lane="2" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25868" lane="6" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25916" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Anna" gender="F" lastname="Cao" nation="GER" license="417196" athleteid="24782">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.73" eventid="5712" heatid="25841" lane="3" />
                <ENTRY entrytime="00:00:51.03" eventid="5728" heatid="25874" lane="2" />
                <ENTRY entrytime="00:01:45.73" eventid="1135" heatid="25896" lane="6" />
                <ENTRY entrytime="00:00:45.23" eventid="5744" heatid="25923" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Anton" gender="M" lastname="Cao" nation="GER" license="417199" athleteid="24787">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.83" eventid="1053" heatid="25749" lane="4" />
                <ENTRY entrytime="00:00:26.68" eventid="5678" heatid="25769" lane="2" />
                <ENTRY entrytime="00:00:30.66" eventid="5694" heatid="25801" lane="5" />
                <ENTRY entrytime="NT" eventid="7701" heatid="25807" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Valentina" gender="F" lastname="Dörner" nation="GER" license="420704" athleteid="25541">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1183" heatid="25814" lane="4" />
                <ENTRY entrytime="NT" eventid="5712" heatid="25833" lane="4" />
                <ENTRY entrytime="NT" eventid="5728" status="DNS" heatid="25864" lane="3" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25887" lane="4" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25913" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Marie" gender="F" lastname="Ehlert" nation="GER" license="382801" athleteid="24792">
              <ENTRIES>
                <ENTRY entrytime="00:03:22.00" eventid="1183" heatid="25818" lane="5" />
                <ENTRY entrytime="00:00:48.73" eventid="5728" heatid="25875" lane="4" />
                <ENTRY entrytime="00:00:36.56" eventid="5744" heatid="25928" lane="1" />
                <ENTRY entrytime="00:00:18.61" eventid="7809" heatid="25955" lane="4" />
                <ENTRY entrytime="00:03:40.00" eventid="5661" heatid="26009" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Tabea" gender="F" lastname="Engelbach" nation="GER" license="419819" athleteid="24798">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25836" lane="5" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25867" lane="4" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25916" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="David" gender="M" lastname="Engler" nation="GER" license="406755" athleteid="24802">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.04" eventid="5702" heatid="25829" lane="5" />
                <ENTRY entrytime="00:00:56.42" eventid="5724" heatid="25857" lane="4" />
                <ENTRY entrytime="00:00:41.00" eventid="5740" heatid="25909" lane="5" />
                <ENTRY entrytime="00:01:55.00" eventid="7773" heatid="25932" lane="3" />
                <ENTRY entrytime="00:00:25.00" eventid="7804" heatid="25949" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Jonas" gender="M" lastname="Erdmann" nation="GER" license="420491" athleteid="24808">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5702" status="DNS" heatid="25821" lane="4" />
                <ENTRY entrytime="NT" eventid="5724" status="DNS" heatid="25852" lane="3" />
                <ENTRY entrytime="NT" eventid="5740" status="DNS" heatid="25898" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Kim" gender="F" lastname="Forster" nation="GER" license="330020" athleteid="24812">
              <ENTRIES>
                <ENTRY entrytime="00:03:05.67" eventid="1183" heatid="25819" lane="6" />
                <ENTRY entrytime="00:00:45.53" eventid="5712" heatid="25847" lane="6" />
                <ENTRY entrytime="00:00:41.19" eventid="5728" heatid="25877" lane="3" />
                <ENTRY entrytime="00:00:48.65" eventid="1123" heatid="25964" lane="3" />
                <ENTRY entrytime="00:01:34.17" eventid="1171" heatid="25979" lane="5" />
                <ENTRY entrytime="00:03:30.46" eventid="5661" heatid="26010" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Viktor" gender="M" lastname="Grin" nation="GER" license="417201" athleteid="24819">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.43" eventid="5702" heatid="25829" lane="1" />
                <ENTRY entrytime="00:00:56.32" eventid="5724" heatid="25858" lane="6" />
                <ENTRY entrytime="00:01:45.67" eventid="1141" heatid="25884" lane="2" />
                <ENTRY entrytime="00:00:45.67" eventid="5740" heatid="25906" lane="3" />
                <ENTRY entrytime="00:01:59.43" eventid="7773" heatid="25932" lane="1" />
                <ENTRY entrytime="00:00:58.93" eventid="1117" heatid="25957" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Rojan" gender="M" lastname="Günes" nation="GER" license="420709" athleteid="25547">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5702" heatid="25821" lane="2" />
                <ENTRY entrytime="NT" eventid="5724" heatid="25853" lane="5" />
                <ENTRY entrytime="NT" eventid="1141" heatid="25878" lane="1" />
                <ENTRY entrytime="NT" eventid="5740" heatid="25899" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Serwan" gender="M" lastname="Günes" nation="GER" license="420706" athleteid="25539">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25745" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Julian" gender="M" lastname="Hampel" nation="GER" license="401463" athleteid="24826">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.56" eventid="5702" heatid="25825" lane="2" />
                <ENTRY entrytime="00:00:51.00" eventid="5724" heatid="25860" lane="4" />
                <ENTRY entrytime="00:00:47.00" eventid="5740" heatid="25906" lane="1" />
                <ENTRY entrytime="00:02:10.00" eventid="7773" heatid="25931" lane="1" />
                <ENTRY entrytime="00:01:05.00" eventid="1117" heatid="25956" lane="3" />
                <ENTRY entrytime="00:01:56.59" eventid="1189" status="DNS" heatid="25984" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Konstantin" gender="M" lastname="Heiden" nation="GER" license="0" athleteid="24833">
              <ENTRIES>
                <ENTRY entrytime="00:00:42.28" eventid="1053" heatid="25747" lane="1" />
                <ENTRY entrytime="00:00:44.05" eventid="5678" heatid="25767" lane="4" />
                <ENTRY entrytime="00:00:42.08" eventid="7691" heatid="25778" lane="2" />
                <ENTRY entrytime="00:00:42.38" eventid="5686" heatid="25791" lane="5" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25798" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Sandra" gender="F" lastname="Herrler" nation="GER" license="414205" athleteid="24839">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.00" eventid="1135" heatid="25891" lane="1" />
                <ENTRY entrytime="00:01:48.00" eventid="7788" heatid="25942" lane="2" />
                <ENTRY entrytime="00:00:57.00" eventid="1123" heatid="25963" lane="6" />
                <ENTRY entrytime="00:02:01.03" eventid="1171" heatid="25976" lane="6" />
                <ENTRY entrytime="00:01:46.81" eventid="1195" heatid="25999" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Hanna" gender="F" lastname="Holtmannspötter" nation="GER" athleteid="25088">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.00" eventid="5712" heatid="25834" lane="3" />
                <ENTRY entrytime="00:01:10.00" eventid="5728" heatid="25866" lane="4" />
                <ENTRY entrytime="00:01:05.00" eventid="5744" heatid="25915" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Hanna" gender="F" lastname="Jonas" nation="GER" license="420708" athleteid="25552">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25833" lane="2" />
                <ENTRY entrytime="NT" eventid="5728" status="DNS" heatid="25864" lane="1" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25887" lane="2" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25912" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Katharina" gender="F" lastname="Kartucha" nation="GER" license="330019" athleteid="24845">
              <ENTRIES>
                <ENTRY entrytime="00:03:59.00" eventid="1183" heatid="25816" lane="5" />
                <ENTRY entrytime="00:01:13.96" eventid="5712" heatid="25835" lane="2" />
                <ENTRY entrytime="00:01:27.76" eventid="5728" heatid="25865" lane="5" />
                <ENTRY entrytime="00:01:54.37" eventid="1135" heatid="25893" lane="4" />
                <ENTRY entrytime="00:01:29.44" eventid="5744" heatid="25913" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Saskia" gender="F" lastname="Klein" nation="GER" athleteid="25080">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25836" lane="4" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25868" lane="5" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25917" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Ella" gender="F" lastname="Kleinert" nation="GER" license="412139" athleteid="24851">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.00" eventid="5664" heatid="25755" lane="3" />
                <ENTRY entrytime="00:00:37.00" eventid="5674" heatid="25764" lane="5" />
                <ENTRY entrytime="00:00:31.97" eventid="5682" heatid="25772" lane="3" />
                <ENTRY entrytime="00:00:32.00" eventid="5690" heatid="25796" lane="3" />
                <ENTRY entrytime="00:00:29.22" eventid="5698" heatid="25806" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Jonathan" gender="M" lastname="Koepnick" nation="GER" license="408297" athleteid="24857">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.69" eventid="5702" heatid="25831" lane="5" />
                <ENTRY entrytime="00:01:53.00" eventid="1141" heatid="25882" lane="3" />
                <ENTRY entrytime="00:01:48.00" eventid="7773" heatid="25933" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="1117" heatid="25957" lane="2" />
                <ENTRY entrytime="00:01:35.00" eventid="1189" heatid="25988" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2005-01-01" firstname="Paul" gender="M" lastname="Kolosowski" nation="GER" license="417223" athleteid="24869">
              <ENTRIES>
                <ENTRY entrytime="00:03:50.32" eventid="1177" heatid="25810" lane="2" />
                <ENTRY entrytime="00:00:56.32" eventid="5702" heatid="25827" lane="4" />
                <ENTRY entrytime="00:00:55.32" eventid="5724" heatid="25858" lane="1" />
                <ENTRY entrytime="00:02:09.09" eventid="1141" heatid="25880" lane="6" />
                <ENTRY entrytime="00:00:59.28" eventid="5740" heatid="25901" lane="3" />
                <ENTRY entrytime="00:01:56.73" eventid="7773" heatid="25932" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Tom" gender="M" lastname="Kossmann" nation="GER" license="0" athleteid="24876">
              <ENTRIES>
                <ENTRY entrytime="00:00:32.34" eventid="1053" heatid="25748" lane="3" />
                <ENTRY entrytime="00:00:34.91" eventid="5678" heatid="25768" lane="3" />
                <ENTRY entrytime="00:00:48.53" eventid="7691" heatid="25777" lane="4" />
                <ENTRY entrytime="00:00:34.81" eventid="5694" heatid="25800" lane="2" />
                <ENTRY entrytime="NT" eventid="7701" heatid="25807" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Ben" gender="M" lastname="Kreibohm" nation="GER" license="0" athleteid="24894">
              <ENTRIES>
                <ENTRY entrytime="00:00:40.41" eventid="5678" heatid="25768" lane="1" />
                <ENTRY entrytime="00:00:44.81" eventid="7691" heatid="25778" lane="6" />
                <ENTRY entrytime="00:00:44.12" eventid="5686" heatid="25791" lane="1" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25797" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Alessia" gender="F" lastname="Köhler" nation="GER" license="399200" athleteid="24863">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.19" eventid="5712" heatid="25845" lane="5" />
                <ENTRY entrytime="00:01:53.00" eventid="1111" heatid="25850" lane="1" />
                <ENTRY entrytime="00:00:36.56" eventid="5744" heatid="25928" lane="6" />
                <ENTRY entrytime="00:00:18.56" eventid="7809" heatid="25955" lane="3" />
                <ENTRY entrytime="00:03:40.00" eventid="5661" heatid="26010" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Madlen" gender="F" lastname="Köthe" nation="GER" license="393115" athleteid="24882">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.84" eventid="5664" heatid="25754" lane="4" />
                <ENTRY entrytime="00:00:24.79" eventid="5682" heatid="25773" lane="5" />
                <ENTRY entrytime="00:00:30.00" eventid="7696" heatid="25785" lane="2" />
                <ENTRY entrytime="00:00:26.09" eventid="5698" heatid="25806" lane="2" />
                <ENTRY entrytime="00:00:34.00" eventid="7706" heatid="25809" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Nina" gender="F" lastname="Köttschau" nation="GER" license="392885" athleteid="24888">
              <ENTRIES>
                <ENTRY entrytime="00:01:55.07" eventid="1135" heatid="25893" lane="5" />
                <ENTRY entrytime="00:01:47.02" eventid="7788" heatid="25942" lane="3" />
                <ENTRY entrytime="00:00:45.14" eventid="1123" heatid="25965" lane="2" />
                <ENTRY entrytime="00:01:45.64" eventid="1171" heatid="25977" lane="2" />
                <ENTRY entrytime="00:01:32.61" eventid="1195" heatid="26002" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Judith" gender="F" lastname="Lerch" nation="GER" license="392892" athleteid="24899">
              <ENTRIES>
                <ENTRY entrytime="00:01:58.75" eventid="1135" heatid="25892" lane="2" />
                <ENTRY entrytime="00:01:50.00" eventid="7788" heatid="25942" lane="1" />
                <ENTRY entrytime="00:00:49.33" eventid="1123" heatid="25964" lane="2" />
                <ENTRY entrytime="00:01:55.33" eventid="1171" heatid="25976" lane="2" />
                <ENTRY entrytime="00:01:41.17" eventid="1195" heatid="26001" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Suljewic" gender="F" lastname="Lina" nation="GER" license="0" athleteid="24905">
              <ENTRIES>
                <ENTRY entrytime="00:00:36.85" eventid="5664" heatid="25754" lane="1" />
                <ENTRY entrytime="00:00:31.44" eventid="5682" heatid="25773" lane="1" />
                <ENTRY entrytime="00:00:41.03" eventid="7696" heatid="25785" lane="6" />
                <ENTRY entrytime="00:00:35.75" eventid="5698" heatid="25805" lane="4" />
                <ENTRY entrytime="NT" eventid="7706" heatid="25808" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Helena Maricosa" gender="F" lastname="Lohmann" nation="GER" license="420492" athleteid="24911">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5728" heatid="25865" lane="1" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25913" lane="2" />
                <ENTRY entrytime="NT" eventid="7809" heatid="25951" lane="1" />
                <ENTRY entrytime="NT" eventid="1171" heatid="25973" lane="2" />
                <ENTRY entrytime="NT" eventid="1195" heatid="25993" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Johanna" gender="F" lastname="Markus" nation="GER" license="0" athleteid="24917">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5664" heatid="25750" lane="4" />
                <ENTRY entrytime="NT" eventid="5682" heatid="25770" lane="1" />
                <ENTRY entrytime="NT" eventid="5690" heatid="25792" lane="3" />
                <ENTRY entrytime="NT" eventid="5698" heatid="25802" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Paolo" gender="M" lastname="Marzo" nation="GER" athleteid="25092">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.00" eventid="5702" heatid="25822" lane="4" />
                <ENTRY entrytime="00:01:10.00" eventid="5740" heatid="25900" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Sarah" gender="F" lastname="Metz" nation="GER" license="382068" athleteid="24922">
              <ENTRIES>
                <ENTRY entrytime="00:01:38.83" eventid="1135" heatid="25897" lane="1" />
                <ENTRY entrytime="00:01:35.38" eventid="7788" heatid="25945" lane="1" />
                <ENTRY entrytime="00:00:45.60" eventid="1123" heatid="25965" lane="5" />
                <ENTRY entrytime="00:01:38.17" eventid="1171" heatid="25978" lane="3" />
                <ENTRY entrytime="00:01:19.47" eventid="1195" heatid="26005" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Julina" gender="F" lastname="Michel" nation="GER" license="404917" athleteid="24928">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.13" eventid="5712" heatid="25843" lane="1" />
                <ENTRY entrytime="00:00:50.10" eventid="5728" heatid="25874" lane="3" />
                <ENTRY entrytime="00:00:44.09" eventid="5744" heatid="25924" lane="6" />
                <ENTRY entrytime="00:01:51.88" eventid="7788" heatid="25941" lane="2" />
                <ENTRY entrytime="00:00:22.78" eventid="7809" heatid="25955" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Phiene" gender="F" lastname="Obermann" nation="GER" license="420707" athleteid="25557">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25834" lane="6" />
                <ENTRY entrytime="NT" eventid="5728" status="DNS" heatid="25864" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Milana" gender="F" lastname="Oeftering" nation="GER" license="406752" athleteid="24934">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.34" eventid="5712" heatid="25841" lane="2" />
                <ENTRY entrytime="00:01:07.83" eventid="5728" heatid="25866" lane="3" />
                <ENTRY entrytime="00:00:53.70" eventid="5744" heatid="25919" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Sebastian" gender="M" lastname="Pendlebury" nation="GER" license="406824" athleteid="24938">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.63" eventid="5702" heatid="25824" lane="6" />
                <ENTRY entrytime="00:01:10.47" eventid="5724" heatid="25854" lane="5" />
                <ENTRY entrytime="00:00:59.06" eventid="5740" heatid="25902" lane="6" />
                <ENTRY entrytime="00:00:29.00" eventid="7804" heatid="25948" lane="6" />
                <ENTRY entrytime="00:02:10.00" eventid="1189" heatid="25982" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lilli" gender="F" lastname="Pikarski" nation="GER" license="419818" athleteid="24944">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.00" eventid="5712" heatid="25835" lane="3" />
                <ENTRY entrytime="00:01:05.00" eventid="5728" heatid="25868" lane="1" />
                <ENTRY entrytime="00:01:00.00" eventid="5744" heatid="25916" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lia" gender="F" lastname="Puzicha" nation="GER" license="390447" athleteid="24948">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.48" eventid="5712" heatid="25840" lane="1" />
                <ENTRY entrytime="00:00:57.70" eventid="5728" heatid="25871" lane="6" />
                <ENTRY entrytime="00:00:49.59" eventid="5744" heatid="25921" lane="1" />
                <ENTRY entrytime="00:02:10.00" eventid="7788" heatid="25939" lane="5" />
                <ENTRY entrytime="00:00:58.00" eventid="1123" heatid="25962" lane="4" />
                <ENTRY entrytime="00:02:10.00" eventid="1171" heatid="25975" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Anna" gender="F" lastname="Ratay" nation="GER" athleteid="25095">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.00" eventid="5712" heatid="25835" lane="6" />
                <ENTRY entrytime="00:01:10.00" eventid="5728" heatid="25866" lane="5" />
                <ENTRY entrytime="00:01:05.00" eventid="5744" heatid="25915" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Wadim" gender="M" lastname="Reiner" nation="GER" license="415619" athleteid="24955">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1141" heatid="25878" lane="5" />
                <ENTRY entrytime="00:00:58.90" eventid="5740" heatid="25902" lane="1" />
                <ENTRY entrytime="NT" eventid="7773" heatid="25930" lane="5" />
                <ENTRY entrytime="00:02:32.17" eventid="1165" heatid="25968" lane="6" />
                <ENTRY entrytime="00:02:33.87" eventid="1189" heatid="25982" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Adrian" gender="M" lastname="Rohn" nation="GER" license="390446" athleteid="24961">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.27" eventid="5702" heatid="25826" lane="3" />
                <ENTRY entrytime="00:00:46.59" eventid="5724" heatid="25862" lane="2" />
                <ENTRY entrytime="00:00:41.68" eventid="5740" heatid="25908" lane="3" />
                <ENTRY entrytime="00:00:25.62" eventid="7804" heatid="25949" lane="1" />
                <ENTRY entrytime="00:01:50.47" eventid="1165" heatid="25969" lane="3" />
                <ENTRY entrytime="00:04:03.00" eventid="5655" heatid="26006" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Luisa" gender="F" lastname="Rübner" nation="GER" license="420493" athleteid="24968">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.12" eventid="5712" heatid="25836" lane="3" />
                <ENTRY entrytime="00:01:01.06" eventid="5728" heatid="25870" lane="1" />
                <ENTRY entrytime="00:00:50.04" eventid="5744" heatid="25920" lane="3" />
                <ENTRY entrytime="00:01:59.54" eventid="7788" heatid="25940" lane="2" />
                <ENTRY entrytime="00:01:59.24" eventid="1195" heatid="25997" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Michael" gender="M" lastname="Rübner" nation="GER" license="385452" athleteid="24974">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.79" eventid="5724" heatid="25857" lane="6" />
                <ENTRY entrytime="00:00:48.73" eventid="5740" heatid="25904" lane="2" />
                <ENTRY entrytime="00:01:58.87" eventid="7773" heatid="25932" lane="5" />
                <ENTRY entrytime="00:00:59.58" eventid="1117" heatid="25957" lane="4" />
                <ENTRY entrytime="00:01:52.66" eventid="1189" heatid="25985" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Massimo" gender="M" lastname="Sauter" nation="GER" license="392205" athleteid="24980">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.00" eventid="5702" heatid="25823" lane="4" />
                <ENTRY entrytime="00:00:55.00" eventid="5724" heatid="25858" lane="2" />
                <ENTRY entrytime="00:00:48.00" eventid="5740" heatid="25905" lane="1" />
                <ENTRY entrytime="00:00:28.00" eventid="7804" heatid="25948" lane="2" />
                <ENTRY entrytime="00:02:00.34" eventid="1189" heatid="25983" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Brian" gender="M" lastname="Schneidt" nation="GER" license="374870" athleteid="24986">
              <ENTRIES>
                <ENTRY entrytime="00:03:14.13" eventid="1177" heatid="25812" lane="6" />
                <ENTRY entrytime="00:00:41.72" eventid="5724" heatid="25863" lane="5" />
                <ENTRY entrytime="00:00:38.70" eventid="5740" heatid="25910" lane="5" />
                <ENTRY entrytime="00:00:20.13" eventid="7804" heatid="25950" lane="2" />
                <ENTRY entrytime="00:03:40.00" eventid="5655" heatid="26007" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Lisa-Joye" gender="F" lastname="Schopf" nation="GER" license="404732" athleteid="24992">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.38" eventid="5712" heatid="25841" lane="5" />
                <ENTRY entrytime="00:00:53.85" eventid="5728" heatid="25873" lane="6" />
                <ENTRY entrytime="00:00:49.19" eventid="5744" heatid="25921" lane="4" />
                <ENTRY entrytime="00:00:26.00" eventid="7809" heatid="25953" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1171" heatid="25976" lane="5" />
                <ENTRY entrytime="00:01:58.00" eventid="1195" heatid="25997" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Leanora" gender="F" lastname="Sebeld" nation="GER" license="414884" athleteid="24999">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.08" eventid="5728" heatid="25872" lane="6" />
                <ENTRY entrytime="00:00:55.10" eventid="5744" heatid="25918" lane="3" />
                <ENTRY entrytime="00:02:05.00" eventid="7788" heatid="25939" lane="2" />
                <ENTRY entrytime="00:00:24.00" eventid="7809" heatid="25954" lane="4" />
                <ENTRY entrytime="00:02:08.00" eventid="1171" heatid="25975" lane="2" />
                <ENTRY entrytime="00:02:05.00" eventid="1195" heatid="25996" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2012-01-01" firstname="Benjamin" gender="M" lastname="Seeger" nation="GER" license="0" athleteid="25006">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1053" heatid="25744" lane="3" />
                <ENTRY entrytime="NT" eventid="5678" heatid="25765" lane="4" />
                <ENTRY entrytime="NT" eventid="5686" heatid="25788" lane="6" />
                <ENTRY entrytime="NT" eventid="5694" heatid="25798" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Veit-Josef" gender="M" lastname="Seidel" nation="GER" license="393117" athleteid="25011">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.00" eventid="5702" heatid="25829" lane="2" />
                <ENTRY entrytime="00:00:53.95" eventid="5724" heatid="25859" lane="2" />
                <ENTRY entrytime="00:00:46.94" eventid="5740" heatid="25906" lane="2" />
                <ENTRY entrytime="00:02:08.00" eventid="7773" heatid="25931" lane="2" />
                <ENTRY entrytime="00:00:26.00" eventid="7804" heatid="25948" lane="4" />
                <ENTRY entrytime="00:01:53.28" eventid="1189" heatid="25985" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Franziska" gender="F" lastname="Selesi" nation="GER" license="0" athleteid="25018">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5682" heatid="25770" lane="2" />
                <ENTRY entrytime="NT" eventid="7696" heatid="25781" lane="3" />
                <ENTRY entrytime="NT" eventid="7706" status="DNS" heatid="25809" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Elisabeth" gender="F" lastname="Strecker" nation="GER" license="406754" athleteid="25022">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.47" eventid="5712" heatid="25840" lane="5" />
                <ENTRY entrytime="00:00:47.59" eventid="5728" heatid="25876" lane="2" />
                <ENTRY entrytime="00:00:46.91" eventid="5744" heatid="25922" lane="2" />
                <ENTRY entrytime="00:01:55.00" eventid="7788" heatid="25941" lane="1" />
                <ENTRY entrytime="00:00:25.00" eventid="7809" heatid="25954" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Mark" gender="M" lastname="Sukhov" nation="GER" license="406821" athleteid="25028">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.75" eventid="5702" heatid="25826" lane="5" />
                <ENTRY entrytime="00:00:51.78" eventid="5724" heatid="25860" lane="5" />
                <ENTRY entrytime="00:00:42.00" eventid="5740" heatid="25908" lane="1" />
                <ENTRY entrytime="00:02:03.00" eventid="7773" heatid="25931" lane="3" />
                <ENTRY entrytime="00:01:03.00" eventid="1117" heatid="25957" lane="5" />
                <ENTRY entrytime="00:01:43.00" eventid="1189" heatid="25986" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Robin" gender="M" lastname="Tiede" nation="GER" license="404730" athleteid="25035">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.93" eventid="1053" heatid="25749" lane="5" />
                <ENTRY entrytime="00:00:30.23" eventid="5678" heatid="25769" lane="1" />
                <ENTRY entrytime="00:00:35.00" eventid="5686" heatid="25791" lane="3" />
                <ENTRY entrytime="00:00:28.44" eventid="5694" heatid="25801" lane="4" />
                <ENTRY entrytime="00:00:28.00" eventid="7701" heatid="25807" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Tobias" gender="M" lastname="Tolba" nation="GER" license="404733" athleteid="25041">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="5702" heatid="25824" lane="5" />
                <ENTRY entrytime="00:00:58.38" eventid="5724" heatid="25857" lane="1" />
                <ENTRY entrytime="00:00:54.97" eventid="5740" heatid="25902" lane="3" />
                <ENTRY entrytime="00:00:26.00" eventid="7804" heatid="25949" lane="6" />
                <ENTRY entrytime="00:02:10.00" eventid="1165" heatid="25968" lane="5" />
                <ENTRY entrytime="00:02:04.72" eventid="1189" heatid="25983" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Laura" gender="F" lastname="Viva" nation="GER" license="420705" athleteid="25560">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5712" heatid="25834" lane="5" />
                <ENTRY entrytime="NT" eventid="1135" heatid="25888" lane="5" />
                <ENTRY entrytime="NT" eventid="5744" heatid="25913" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Adrian" gender="M" lastname="Vorrat" nation="GER" license="392206" athleteid="25048">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.00" eventid="5702" heatid="25826" lane="6" />
                <ENTRY entrytime="00:00:50.00" eventid="5724" heatid="25861" lane="2" />
                <ENTRY entrytime="00:00:48.00" eventid="5740" heatid="25905" lane="5" />
                <ENTRY entrytime="00:00:26.00" eventid="7804" heatid="25948" lane="3" />
                <ENTRY entrytime="00:02:02.50" eventid="1165" heatid="25968" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Malin" gender="F" lastname="Wachter" nation="GER" license="393237" athleteid="25054">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.34" eventid="5712" status="DNS" heatid="25846" lane="6" />
                <ENTRY entrytime="00:00:44.00" eventid="5728" status="DNS" heatid="25877" lane="5" />
                <ENTRY entrytime="00:00:36.67" eventid="5744" status="DNS" heatid="25927" lane="4" />
                <ENTRY entrytime="00:00:19.64" eventid="7809" status="DNS" heatid="25955" lane="2" />
                <ENTRY entrytime="00:01:53.29" eventid="1171" status="DNS" heatid="25977" lane="6" />
                <ENTRY entrytime="00:03:40.00" eventid="5661" status="DNS" heatid="26010" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Mara Malin" gender="F" lastname="Walther" nation="GER" license="362627" athleteid="25061">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.94" eventid="5712" heatid="25844" lane="2" />
                <ENTRY entrytime="00:00:52.16" eventid="5728" heatid="25873" lane="4" />
                <ENTRY entrytime="00:00:45.70" eventid="5744" heatid="25923" lane="2" />
                <ENTRY entrytime="00:01:00.06" eventid="1123" heatid="25962" lane="5" />
                <ENTRY entrytime="00:04:15.00" eventid="5661" heatid="26008" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Sophia" gender="F" lastname="Walther" nation="GER" license="414879" athleteid="25067">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.22" eventid="5712" heatid="25841" lane="4" />
                <ENTRY entrytime="00:01:01.77" eventid="5728" heatid="25869" lane="3" />
                <ENTRY entrytime="00:00:54.88" eventid="5744" heatid="25919" lane="1" />
                <ENTRY entrytime="00:00:26.00" eventid="7809" heatid="25953" lane="2" />
                <ENTRY entrytime="00:02:08.00" eventid="1195" heatid="25996" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Helena" gender="F" lastname="Willared" nation="GER" license="368438" athleteid="25073">
              <ENTRIES>
                <ENTRY entrytime="00:01:54.42" eventid="1135" heatid="25893" lane="2" />
                <ENTRY entrytime="00:01:45.47" eventid="7788" heatid="25943" lane="5" />
                <ENTRY entrytime="00:00:49.44" eventid="1123" heatid="25964" lane="5" />
                <ENTRY entrytime="00:01:44.27" eventid="1171" heatid="25977" lane="4" />
                <ENTRY entrytime="00:01:32.74" eventid="1195" heatid="26002" lane="1" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="8" agetotalmax="-1" agetotalmin="-1" gender="X">
              <ENTRIES>
                <ENTRY entrytime="00:01:47.65" eventid="23774" heatid="25946" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="24986" number="1" />
                    <RELAYPOSITION athleteid="24741" number="2" />
                    <RELAYPOSITION athleteid="24863" number="3" />
                    <RELAYPOSITION athleteid="24792" number="4" />
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
          <OFFICIALS>
            <OFFICIAL officialid="17182" firstname="Claudia" gender="F" lastname="Bachmann" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26028" firstname="Peter" gender="M" lastname="Baumann" nation="GER">
              <CONTACT city="SV Franken" />
            </OFFICIAL>
            <OFFICIAL officialid="26043" firstname="Julian" gender="M" lastname="Beyer" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26115" firstname="Kristin" gender="F" lastname="Braun-Klimpel" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23617" firstname="Andreas" gender="M" lastname="Distler" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="17202" firstname="Frank" gender="M" lastname="Emmerlich" nation="GER" />
            <OFFICIAL officialid="26101" firstname="Donald" gender="M" lastname="Forster" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23656" firstname="Torsten" gender="M" lastname="Heiden" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23601" firstname="Ralph" gender="M" lastname="Jonscher" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="17220" firstname="Nicole" gender="F" lastname="Kleinhenz" nation="GER" />
            <OFFICIAL officialid="26103" firstname="Eva-Katharina" gender="F" lastname="Krämer" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23603" firstname="Roland" gender="M" lastname="Köhler" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26058" firstname="Sedat" gender="M" lastname="Köthe" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="17210" firstname="Sadet" gender="F" lastname="Kötne" nation="GER" />
            <OFFICIAL officialid="26095" firstname="Wibke" gender="F" lastname="Lerch" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23678" firstname="Matthias" gender="M" lastname="Meixner" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26055" firstname="Julian" gender="M" lastname="Messel" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26066" firstname="Katharina" gender="F" lastname="Roth" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23613" firstname="Nils" gender="M" lastname="Rudolph" nation="GER">
              <CONTACT city="TB Erlangen" />
            </OFFICIAL>
            <OFFICIAL officialid="17221" firstname="Sabine" gender="F" lastname="Sandner-Dewdney" nation="GER" />
            <OFFICIAL officialid="17211" firstname="Ulrike" gender="F" lastname="Schall" nation="GER" />
            <OFFICIAL officialid="17180" firstname="Ulrike" gender="F" lastname="Scharnweber" nation="GER" />
            <OFFICIAL officialid="17203" firstname="Florian" gender="M" lastname="Schilling" nation="GER" />
            <OFFICIAL officialid="26102" firstname="Claudia" gender="F" lastname="Schopf" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26107" firstname="Justin" gender="F" lastname="Schreiber" nation="GER">
              <CONTACT city="VfL Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="23669" firstname="Jobst" gender="M" lastname="Schuseil" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26034" firstname="Elisabeth" gender="F" lastname="Seilbold" nation="GER">
              <CONTACT city="SV Franken" />
            </OFFICIAL>
            <OFFICIAL officialid="23579" firstname="Sybille" gender="F" lastname="Streicher" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="17213" firstname="Mike" gender="M" lastname="Sturm" nation="GER" />
            <OFFICIAL officialid="23615" firstname="Xenia" gender="F" lastname="Sukhof" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="26051" firstname="Joachim" gender="M" lastname="Suljewic" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23676" firstname="Joachim" gender="M" lastname="Suljewic" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23769" firstname="Birgit" gender="F" lastname="Thiele" nation="GER">
              <CONTACT city="TSV 1846 Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="17222" firstname="Larissa" gender="F" lastname="Tillner" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="23657" firstname="Timo" gender="M" lastname="Wasmuth" nation="GER">
              <CONTACT city="TSV Altenfurt" />
            </OFFICIAL>
            <OFFICIAL officialid="26118" firstname="Anja" gender="F" lastname="Willard" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
            <OFFICIAL officialid="17206" firstname="Petra" gender="F" lastname="Wormser" nation="GER">
              <CONTACT city="SG Mittelfranken" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="5541" nation="GER" region="02" clubid="7909" name="SG Nordoberpfalz" />
        <CLUB type="CLUB" code="4305" nation="GER" region="02" clubid="7958" name="SG Oberland Penzberg" />
        <CLUB type="CLUB" code="6621" nation="GER" region="02" clubid="7924" name="SG Rödental" />
        <CLUB type="CLUB" code="6423" nation="GER" region="02" clubid="7931" name="SG Stadtwerke München">
          <OFFICIALS>
            <OFFICIAL officialid="23670" firstname="Karin" gender="F" lastname="Bartel" nation="GER">
              <CONTACT city="SG Stadtwerke München" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4958" nation="GER" region="02" clubid="7944" name="SSG 81 Erlangen">
          <OFFICIALS>
            <OFFICIAL officialid="26116" firstname="Ditmar" gender="M" lastname="Asse" nation="GER">
              <CONTACT city="SSG 81 Erlangen" />
            </OFFICIAL>
            <OFFICIAL officialid="17207" firstname="Roland" gender="M" lastname="Beer" nation="GER" />
            <OFFICIAL officialid="17216" firstname="Katharina" gender="F" lastname="Brem" nation="GER">
              <CONTACT city="SSG Erlangen" />
            </OFFICIAL>
            <OFFICIAL officialid="17219" firstname="Nowak" gender="M" lastname="Götz" nation="GER">
              <CONTACT city="SSG 81 Erlangen" />
            </OFFICIAL>
            <OFFICIAL officialid="23768" firstname="Isabella" gender="F" lastname="Kaufmann" nation="GER">
              <CONTACT city="SSG 81 Erlangen" />
            </OFFICIAL>
            <OFFICIAL officialid="23761" firstname="Manfred" gender="M" lastname="Kreißel" nation="GER">
              <CONTACT city="TB Erlangen" />
            </OFFICIAL>
            <OFFICIAL officialid="23765" firstname="Katrin" gender="F" lastname="Rudolph" nation="GER">
              <CONTACT city="TB Erlangen" />
            </OFFICIAL>
            <OFFICIAL officialid="23764" firstname="Nele" gender="F" lastname="Rudolph" nation="GER">
              <CONTACT city="TB Erlangen" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4328" nation="GER" region="02" clubid="7957" name="SSG Bad Reichenhall im BGL e.V." shortname="SSG Bad Reichenhall im BGL e.V" />
        <CLUB type="CLUB" code="6695" nation="GER" region="02" clubid="7969" name="SSG Coburg" />
        <CLUB type="CLUB" code="4329" nation="GER" region="02" clubid="7929" name="SSG Günzburg-Leipheim" />
        <CLUB type="CLUB" code="4330" nation="GER" region="02" clubid="7922" name="SSG Neptun Germering e.V." />
        <CLUB type="CLUB" code="4331" nation="GER" region="02" clubid="7937" name="SSKC Poseidon Aschaffenburg" />
        <CLUB type="CLUB" code="4332" nation="GER" region="02" clubid="7946" name="SSV Forchheim">
          <OFFICIALS>
            <OFFICIAL officialid="17217" firstname="Denisa" gender="F" lastname="Kisberi" nation="GER">
              <CONTACT city="SSV Forchheim" />
            </OFFICIAL>
            <OFFICIAL officialid="17205" firstname="Lidia" gender="F" lastname="Pira" nation="GER" />
            <OFFICIAL officialid="17186" firstname="Stefan" gender="M" lastname="Wagner" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4336" nation="GER" region="02" clubid="7916" name="SSV Höchstädt" />
        <CLUB type="CLUB" code="4362" nation="GER" region="02" clubid="7890" name="SV 77 Neufahrn" />
        <CLUB type="CLUB" code="4343" nation="GER" region="02" clubid="7927" name="SV Arnbruck" />
        <CLUB type="CLUB" code="4347" nation="GER" region="02" clubid="7918" name="SV Bayreuth" />
        <CLUB type="CLUB" nation="GER" region="02" clubid="25537" name="SV Franken" />
        <CLUB type="CLUB" code="4385" nation="GER" region="02" clubid="7891" name="SV Fürstenfeldbrucker Wasserratten e.V." shortname="SV Fürstenfeldbrucker Wasserra" />
        <CLUB type="CLUB" code="4356" nation="GER" region="02" clubid="7899" name="SV GR.-W. Holzkirchen" />
        <CLUB type="CLUB" code="4357" nation="GER" region="02" clubid="7894" name="SV Grafing-Ebersberg" />
        <CLUB type="CLUB" code="5713" nation="GER" region="02" clubid="7971" name="SV Hengersberg" />
        <CLUB type="CLUB" code="4341" nation="GER" region="02" clubid="7915" name="SV Hof 1911 e. V." />
        <CLUB type="CLUB" code="4360" nation="GER" region="02" clubid="7952" name="SV Lohhof" />
        <CLUB type="CLUB" code="4364" nation="GER" region="02" clubid="7900" name="SV Ottobrunn 1970 e.V." />
        <CLUB type="CLUB" code="4374" nation="GER" region="02" clubid="7943" name="SV Schwabach" />
        <CLUB type="CLUB" code="4384" nation="GER" region="02" clubid="7898" name="SV Wacker Burghausen" />
        <CLUB type="CLUB" code="4387" nation="GER" region="02" clubid="7932" name="SV Weiden" />
        <CLUB type="CLUB" code="4339" nation="GER" region="02" clubid="7960" name="SV Würzburg 05" />
        <CLUB type="CLUB" code="5806" nation="GER" region="02" clubid="7935" name="Team Buron Kaufbeuren" />
        <CLUB type="CLUB" code="4405" nation="GER" region="02" clubid="7897" name="TSG Kleinostheim" />
        <CLUB type="CLUB" code="6655" nation="GER" region="02" clubid="7904" name="TSG Nürnberg">
          <ATHLETES>
            <ATHLETE birthdate="2011-01-01" firstname="Leni" gender="F" lastname="Amadasun" nation="GER" license="0" athleteid="25111">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.00" eventid="5664" heatid="25755" lane="4" />
                <ENTRY entrytime="00:00:30.00" eventid="5674" heatid="25764" lane="3" />
                <ENTRY entrytime="00:00:23.00" eventid="5682" heatid="25773" lane="2" />
                <ENTRY entrytime="00:00:30.00" eventid="7696" heatid="25785" lane="5" />
                <ENTRY entrytime="00:00:26.00" eventid="5698" heatid="25806" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="7706" heatid="25809" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Alexey" gender="M" lastname="Antonkin" nation="GER" license="392619" athleteid="25118">
              <ENTRIES>
                <ENTRY entrytime="00:03:16.33" eventid="1177" heatid="25811" lane="3" />
                <ENTRY entrytime="00:00:56.14" eventid="5702" heatid="25828" lane="6" />
                <ENTRY entrytime="00:02:00.00" eventid="1103" heatid="25848" lane="6" />
                <ENTRY entrytime="00:01:53.92" eventid="1165" heatid="25969" lane="2" />
                <ENTRY entrytime="00:03:54.69" eventid="5655" heatid="26006" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2011-01-01" firstname="Sandrine" gender="F" lastname="Fuchs" nation="GER" license="0" athleteid="25124">
              <ENTRIES>
                <ENTRY entrytime="00:00:37.00" eventid="5674" heatid="25764" lane="2" />
                <ENTRY entrytime="00:00:33.00" eventid="5682" heatid="25772" lane="5" />
                <ENTRY entrytime="00:00:40.00" eventid="7696" heatid="25785" lane="1" />
                <ENTRY entrytime="00:00:37.00" eventid="5698" heatid="25805" lane="5" />
                <ENTRY entrytime="00:00:40.00" eventid="7706" heatid="25809" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-01-01" firstname="Lorena" gender="F" lastname="Graz" nation="GER" license="392620" athleteid="25130">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.91" eventid="5712" heatid="25843" lane="4" />
                <ENTRY entrytime="00:00:51.20" eventid="5728" heatid="25874" lane="5" />
                <ENTRY entrytime="00:00:42.79" eventid="5744" heatid="25924" lane="5" />
                <ENTRY entrytime="00:00:55.28" eventid="1123" heatid="25963" lane="2" />
                <ENTRY entrytime="00:01:46.54" eventid="1195" heatid="25999" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Luis" gender="M" lastname="Heik" nation="GER" license="377052" athleteid="25136">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.64" eventid="5702" heatid="25830" lane="6" />
                <ENTRY entrytime="00:01:54.39" eventid="1141" heatid="25882" lane="6" />
                <ENTRY entrytime="00:01:45.00" eventid="7773" heatid="25933" lane="5" />
                <ENTRY entrytime="00:00:22.00" eventid="7804" heatid="25950" lane="1" />
                <ENTRY entrytime="00:01:42.29" eventid="1189" heatid="25987" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2009-07-06" firstname="Cedrik" gender="M" lastname="Kreik" nation="GER" license="99999" athleteid="26016">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.92" eventid="5702" />
                <ENTRY entrytime="NT" eventid="1103" />
                <ENTRY entrytime="00:01:47.17" eventid="1141" />
                <ENTRY entrytime="00:00:46.17" eventid="1117" />
                <ENTRY entrytime="00:01:32.22" eventid="1189" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Valeria Alexandra" gender="F" lastname="Nekrasov" nation="GER" license="392621" athleteid="25142">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.00" eventid="5712" heatid="25846" lane="1" />
                <ENTRY entrytime="00:01:50.00" eventid="1135" heatid="25894" lane="4" />
                <ENTRY entrytime="00:01:45.00" eventid="7788" heatid="25943" lane="3" />
                <ENTRY entrytime="00:00:50.00" eventid="1123" heatid="25963" lane="3" />
                <ENTRY entrytime="00:01:35.67" eventid="1195" heatid="26001" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Victoria" gender="F" lastname="Nekrasov" nation="GER" license="359482" athleteid="25148">
              <ENTRIES>
                <ENTRY entrytime="00:02:49.85" eventid="1183" heatid="25820" lane="5" />
                <ENTRY entrytime="00:01:26.95" eventid="1111" heatid="25851" lane="2" />
                <ENTRY entrytime="00:01:35.43" eventid="7788" heatid="25945" lane="6" />
                <ENTRY entrytime="00:00:36.48" eventid="1123" heatid="25966" lane="3" />
                <ENTRY entrytime="00:03:07.25" eventid="5661" heatid="26011" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Tobias" gender="M" lastname="Rhau" nation="GER" athleteid="25166">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.00" eventid="5702" status="DNS" heatid="25822" lane="3" />
                <ENTRY entrytime="00:02:20.00" eventid="1141" heatid="25879" lane="4" />
                <ENTRY entrytime="00:01:10.00" eventid="5740" heatid="25900" lane="4" />
                <ENTRY entrytime="00:00:35.00" eventid="7804" status="DNS" heatid="25947" lane="1" />
                <ENTRY entrytime="00:02:15.00" eventid="1189" status="DNS" heatid="25982" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-01-01" firstname="Lena" gender="F" lastname="Schreiber" nation="GER" license="392618" athleteid="25154">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.20" eventid="5712" heatid="25840" lane="2" />
                <ENTRY entrytime="00:02:00.00" eventid="1135" heatid="25892" lane="1" />
                <ENTRY entrytime="00:02:15.00" eventid="7788" heatid="25938" lane="3" />
                <ENTRY entrytime="00:00:35.00" eventid="7809" heatid="25952" lane="5" />
                <ENTRY entrytime="00:02:00.00" eventid="1195" heatid="25997" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Jakob" gender="M" lastname="Sickmüller" nation="GER" license="359484" athleteid="25160">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.00" eventid="5702" heatid="25831" lane="2" />
                <ENTRY entrytime="00:00:50.00" eventid="5724" heatid="25861" lane="5" />
                <ENTRY entrytime="00:00:44.76" eventid="5740" heatid="25907" lane="2" />
                <ENTRY entrytime="00:00:22.00" eventid="7804" heatid="25950" lane="5" />
                <ENTRY entrytime="00:01:50.00" eventid="1189" heatid="25985" lane="4" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="26104" firstname="Mikhail" gender="M" lastname="Antonkin" nation="GER">
              <CONTACT city="TSG Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="26053" firstname="Carry" gender="F" lastname="Fuchs" nation="GER">
              <CONTACT city="TSG Nürnberg" />
            </OFFICIAL>
            <OFFICIAL officialid="17179" firstname="Antonkin" gender="M" lastname="Mikhail" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4407" nation="GER" region="02" clubid="7920" name="TSG Stadtbergen 1892" />
        <CLUB type="CLUB" code="4439" nation="GER" region="02" clubid="7910" name="TSV - Eintracht Karlsfeld" />
        <CLUB type="CLUB" code="4411" nation="GER" region="02" clubid="7884" name="TSV 1847 Weilheim" />
        <CLUB type="CLUB" code="4412" nation="GER" region="02" clubid="7948" name="TSV 1860 Ansbach">
          <OFFICIALS>
            <OFFICIAL officialid="23612" firstname="Steffi" gender="M" lastname="Konrath" nation="GER">
              <CONTACT city="TSV Ansbach" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4413" nation="GER" region="02" clubid="7901" name="TSV 1860 Rosenheim" />
        <CLUB type="CLUB" code="5075" nation="GER" region="02" clubid="7885" name="TSV 1862 Bad Reichenhall" />
        <CLUB type="CLUB" code="4417" nation="GER" region="02" clubid="7887" name="TSV 1862 Friedberg" />
        <CLUB type="CLUB" code="4421" nation="GER" region="02" clubid="7938" name="TSV 1863 Marktoberdorf" />
        <CLUB type="CLUB" code="4445" nation="GER" region="02" clubid="7936" name="TSV 1909 Gersthofen" />
        <CLUB type="CLUB" code="5460" nation="GER" region="02" clubid="7939" name="TSV Delphine Abensberg" />
        <CLUB type="CLUB" code="4441" nation="GER" region="02" clubid="7956" name="TSV Erding" />
        <CLUB type="CLUB" code="4513" nation="GER" region="02" clubid="7895" name="TSV Haar" />
        <CLUB type="CLUB" code="4452" nation="GER" region="02" clubid="7905" name="TSV Hohenbrunn-Riemerl.">
          <OFFICIALS>
            <OFFICIAL officialid="23578" firstname="Claudia" gender="M" lastname="Hermeking" nation="GER">
              <CONTACT city="TSV Hohenbrunn-Riem" />
            </OFFICIAL>
            <OFFICIAL officialid="23590" firstname="Kathi" gender="F" lastname="Schweiger" nation="GER">
              <CONTACT city="TSV Hohenbrunn-Riem" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="6628" nation="GER" region="02" clubid="7893" name="TSV Indersdorf 1907 e.V." />
        <CLUB type="CLUB" code="4415" nation="GER" region="02" clubid="7925" name="TSV Mindelheim" />
        <CLUB type="CLUB" code="4420" nation="GER" region="02" clubid="7941" name="TSV Neuburg" />
        <CLUB type="CLUB" code="4484" nation="GER" region="02" clubid="7928" name="TSV Schwabmünchen" />
        <CLUB type="CLUB" code="4488" nation="GER" region="02" clubid="7888" name="TSV Solln" />
        <CLUB type="CLUB" code="6408" nation="GER" region="02" clubid="7949" name="TSV Stein">
          <OFFICIALS>
            <OFFICIAL officialid="17174" firstname="Tobias" gender="M" lastname="Kloth" nation="GER">
              <CONTACT city="TSV" />
            </OFFICIAL>
            <OFFICIAL officialid="17184" firstname="Andreas" gender="M" lastname="Mittmann" nation="GER" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4492" nation="GER" region="02" clubid="7889" name="TSV Vaterstetten" />
        <CLUB type="CLUB" code="4502" nation="GER" region="02" clubid="7903" name="TSV Zirndorf">
          <ATHLETES>
            <ATHLETE birthdate="2005-01-01" firstname="Jana" gender="F" lastname="Ammon" nation="GER" license="398728" athleteid="23839">
              <ENTRIES>
                <ENTRY entrytime="00:03:25.00" eventid="1183" status="DNS" heatid="25817" lane="4" />
                <ENTRY entrytime="00:00:52.94" eventid="5712" status="DNS" heatid="25844" lane="6" />
                <ENTRY entrytime="00:00:51.59" eventid="5728" status="DNS" heatid="25874" lane="6" />
                <ENTRY entrytime="00:00:41.63" eventid="5744" status="DNS" heatid="25925" lane="1" />
                <ENTRY entrytime="00:01:51.50" eventid="1195" status="DNS" heatid="25998" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Marco" gender="M" lastname="Ammon" nation="GER" license="398727" athleteid="23845">
              <ENTRIES>
                <ENTRY entrytime="00:01:58.94" eventid="1141" heatid="25881" lane="5" />
                <ENTRY entrytime="00:00:43.50" eventid="5740" heatid="25907" lane="3" />
                <ENTRY entrytime="00:01:45.00" eventid="7773" heatid="25933" lane="4" />
                <ENTRY entrytime="00:00:48.25" eventid="1117" heatid="25959" lane="5" />
                <ENTRY entrytime="00:01:35.09" eventid="1189" heatid="25988" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Veit" gender="M" lastname="Bestle" nation="GER" license="398730" athleteid="23851">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.68" eventid="5702" heatid="25831" lane="6" />
                <ENTRY entrytime="00:00:54.50" eventid="5724" heatid="25858" lane="3" />
                <ENTRY entrytime="00:01:55.97" eventid="1141" heatid="25881" lane="3" />
                <ENTRY entrytime="00:00:41.44" eventid="5740" heatid="25909" lane="1" />
                <ENTRY entrytime="00:01:39.62" eventid="1189" heatid="25988" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2008-01-01" firstname="Amélie Marianne" gender="F" lastname="Blumenthal Haz" nation="GER" license="403953" athleteid="23857">
              <ENTRIES>
                <ENTRY entrytime="00:03:25.00" eventid="1183" heatid="25817" lane="3" />
                <ENTRY entrytime="00:01:55.50" eventid="1111" heatid="25849" lane="3" />
                <ENTRY entrytime="00:01:47.94" eventid="7788" heatid="25942" lane="4" />
                <ENTRY entrytime="00:00:22.00" eventid="7809" heatid="25955" lane="5" />
                <ENTRY entrytime="00:01:35.13" eventid="1195" heatid="26001" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2010-10-27" firstname="Mia" gender="F" lastname="Großhauser" nation="GER" license="420483" athleteid="23838">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.00" eventid="5712" heatid="25839" lane="5" />
                <ENTRY entrytime="00:02:21.60" eventid="1135" heatid="25889" lane="6" />
                <ENTRY entrytime="00:00:55.00" eventid="5744" heatid="25919" lane="6" />
                <ENTRY entrytime="00:02:05.00" eventid="1195" heatid="25996" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Jana" gender="F" lastname="Gömmel" nation="GER" license="355570" athleteid="23863">
              <ENTRIES>
                <ENTRY entrytime="00:03:00.00" eventid="1183" heatid="25819" lane="2" />
                <ENTRY entrytime="00:00:45.00" eventid="5728" heatid="25877" lane="6" />
                <ENTRY entrytime="00:00:37.00" eventid="5744" heatid="25927" lane="5" />
                <ENTRY entrytime="00:01:42.37" eventid="7788" status="DNS" heatid="25944" lane="5" />
                <ENTRY entrytime="00:01:20.00" eventid="1195" heatid="26004" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Tim" gender="M" lastname="Krauß" nation="GER" license="407216" athleteid="23875">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.69" eventid="5702" heatid="25826" lane="4" />
                <ENTRY entrytime="00:01:04.37" eventid="5724" heatid="25855" lane="1" />
                <ENTRY entrytime="00:02:00.00" eventid="1141" heatid="25880" lane="3" />
                <ENTRY entrytime="00:00:57.94" eventid="5740" heatid="25902" lane="4" />
                <ENTRY entrytime="00:01:55.00" eventid="1189" heatid="25985" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2007-01-01" firstname="Josefine" gender="F" lastname="Mendler" nation="GER" license="420484" athleteid="24058">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.60" eventid="1195" heatid="25995" lane="2" />
                <ENTRY entrytime="00:01:08.10" eventid="5712" heatid="25837" lane="6" />
                <ENTRY entrytime="00:02:21.60" eventid="1135" heatid="25889" lane="1" />
                <ENTRY entrytime="00:01:02.42" eventid="5744" heatid="25916" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Simona" gender="F" lastname="Paschold" nation="GER" license="398731" athleteid="23881">
              <ENTRIES>
                <ENTRY entrytime="00:03:00.00" eventid="1183" heatid="25819" lane="4" />
                <ENTRY entrytime="00:00:45.16" eventid="5712" heatid="25847" lane="1" />
                <ENTRY entrytime="00:01:42.53" eventid="1135" heatid="25896" lane="4" />
                <ENTRY entrytime="00:00:35.47" eventid="5744" heatid="25928" lane="5" />
                <ENTRY entrytime="00:01:22.57" eventid="1195" heatid="26004" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE birthdate="2006-01-01" firstname="Yannis" gender="M" lastname="Spath" nation="GER" license="385212" athleteid="23887">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.34" eventid="5702" heatid="25830" lane="1" />
                <ENTRY entrytime="00:00:55.00" eventid="5724" heatid="25858" lane="4" />
                <ENTRY entrytime="00:00:40.52" eventid="5740" heatid="25909" lane="4" />
                <ENTRY entrytime="00:01:49.04" eventid="7773" heatid="25933" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="26110" firstname="Wolfgang" gender="M" lastname="Ammon" nation="GER">
              <CONTACT city="TSV Zirndorf" />
            </OFFICIAL>
            <OFFICIAL officialid="26106" firstname="Ngela" gender="F" lastname="Gömmel" nation="GER">
              <CONTACT city="TSV Zirndorf" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="4529" nation="GER" region="02" clubid="7933" name="Turnverein Münchberg" />
        <CLUB type="CLUB" code="5107" nation="GER" region="02" clubid="7963" name="TV 1860 Immenstadt" />
        <CLUB type="CLUB" code="4530" nation="GER" region="02" clubid="7964" name="TV 1862 Passau" />
        <CLUB type="CLUB" code="6812" nation="GER" region="02" clubid="7921" name="TV Kempten" />
        <CLUB type="CLUB" code="4562" nation="GER" region="02" clubid="7906" name="TV Parsberg" />
        <CLUB type="CLUB" code="4523" nation="GER" region="02" clubid="7926" name="TV-Lindenberg" />
        <CLUB type="CLUB" code="4593" nation="GER" region="02" clubid="7968" name="VfL 1860 Spfr. Bad Neustadt" />
        <CLUB type="CLUB" code="4598" nation="GER" region="02" clubid="7934" name="VfL Piranhas Waldkraiburg" />
        <CLUB type="CLUB" code="4595" nation="GER" region="02" clubid="7913" name="VFL-Kaufering" />
        <CLUB type="CLUB" code="4639" nation="GER" region="02" clubid="7955" name="WSV Bad Tölz">
          <OFFICIALS>
            <OFFICIAL officialid="23766" firstname="Maria" gender="F" lastname="Vollmer" nation="GER">
              <CONTACT city="WSV Bad Tölz" />
            </OFFICIAL>
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
